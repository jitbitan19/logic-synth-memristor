// Benchmark "./input/c7552" written by ABC on Thu Aug  8 02:45:58 2024

module c7552  ( 
    G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47,
    G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65,
    G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83,
    G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110,
    G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, G133, G134,
    G135, G138, G141, G144, G147, G150, G151, G152, G153, G154, G155, G156,
    G157, G158, G159, G160, G161, G162, G163, G164, G165, G166, G167, G168,
    G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, G179, G180,
    G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G216,
    G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, G227, G228,
    G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, G239, G240,
    G339, G1197, G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496,
    G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253,
    G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743,
    G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432,
    G4437, G4526, G4528,
    G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399  );
  input  G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41,
    G44, G47, G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63,
    G64, G65, G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81,
    G82, G83, G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106,
    G109, G110, G111, G112, G113, G114, G115, G118, G121, G124, G127, G130,
    G133, G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154,
    G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165, G166,
    G167, G168, G169, G170, G171, G172, G173, G174, G175, G176, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G187, G188, G189, G190,
    G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202,
    G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214,
    G215, G216, G217, G218, G219, G220, G221, G222, G223, G224, G225, G226,
    G227, G228, G229, G230, G231, G232, G233, G234, G235, G236, G237, G238,
    G239, G240, G339, G1197, G1455, G1459, G1462, G1469, G1480, G1486,
    G1492, G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239,
    G2247, G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729,
    G3737, G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420,
    G4427, G4432, G4437, G4526, G4528;
  output G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399;
  wire new_G400_, new_G1184_, new_G1501_, new_G2857_, new_G4442_, new_G4514_,
    new_G401_, new_G573_, new_G574_, new_G575_, new_G1178_, new_G1186_,
    new_G1192_, new_G1198_, new_G1205_, new_G1206_, new_G1207_, new_G1210_,
    new_G1458_, new_G1461_, new_G1464_, new_G1471_, new_G1475_, new_G1482_,
    new_G1488_, new_G1495_, new_G1499_, new_G1500_, new_G1503_, new_G1512_,
    new_G1518_, new_G1524_, new_G1535_, new_G1541_, new_G2207_, new_G2210_,
    new_G2213_, new_G2220_, new_G2226_, new_G2232_, new_G2238_, new_G2241_,
    new_G2249_, new_G2255_, new_G2258_, new_G2828_, new_G3700_, new_G3703_,
    new_G3707_, new_G3713_, new_G3719_, new_G3725_, new_G3731_, new_G3739_,
    new_G3745_, new_G3751_, new_G4121_, new_G4396_, new_G4402_, new_G4407_,
    new_G4412_, new_G4417_, new_G4422_, new_G4429_, new_G4434_, new_G4439_,
    new_G4833_, new_G2876_, new_G2878_, new_G1519_, new_G2871_, new_G2883_,
    new_G280_, new_G4839_, new_G572_, new_G581_, new_G587_, new_G601_,
    new_G606_, new_G650_, new_G657_, new_G671_, new_G678_, new_G777_,
    new_G1115_, new_G1336_, new_G1350_, new_G1477_, new_G1507_, new_G1514_,
    new_G1530_, new_G2259_, new_G2833_, new_G2872_, new_G2886_, new_G2892_,
    new_G2905_, new_G2909_, new_G3622_, new_G3635_, new_G3755_, new_G4640_,
    new_G4653_, new_G4873_, new_G4876_, new_G4881_, new_G4889_, new_G4905_,
    new_G4916_, new_G4921_, new_G5175_, new_G5178_, new_G5186_, new_G5191_,
    new_G5199_, new_G5215_, new_G5223_, new_G5393_, new_G5401_, new_G5409_,
    new_G5417_, new_G5425_, new_G5433_, new_G5441_, new_G5449_, new_G5457_,
    new_G5745_, new_G5753_, new_G5761_, new_G5769_, new_G5777_, new_G5785_,
    new_G5793_, new_G5801_, new_G5809_, new_G5865_, new_G5873_, new_G5881_,
    new_G5889_, new_G5897_, new_G5905_, new_G5913_, new_G5921_, new_G5985_,
    new_G5993_, new_G6001_, new_G6009_, new_G6017_, new_G6025_, new_G6033_,
    new_G6041_, new_G6514_, new_G6554_, new_G6567_, new_G6575_, new_G6583_,
    new_G6591_, new_G6599_, new_G6607_, new_G6615_, new_G6623_, new_G6631_,
    new_G6853_, new_G6861_, new_G6869_, new_G6877_, new_G6885_, new_G6893_,
    new_G6901_, new_G6909_, new_G6917_, new_G784_, new_G1014_, new_G3221_,
    new_G4913_, new_G4929_, new_G5183_, new_G5231_, new_G6511_, new_G615_,
    new_G594_, new_G611_, new_G617_, new_G619_, new_G621_, new_G623_,
    new_G625_, new_G627_, new_G664_, new_G685_, new_G691_, new_G693_,
    new_G695_, new_G697_, new_G699_, new_G701_, new_G703_, new_G705_,
    new_G707_, new_G709_, new_G4879_, new_G4880_, new_G4887_, new_G4895_,
    new_G4911_, new_G4920_, new_G4927_, new_G5181_, new_G5182_, new_G5190_,
    new_G5197_, new_G5205_, new_G5221_, new_G5229_, new_G1343_, new_G1357_,
    new_G1364_, new_G1366_, new_G1368_, new_G1370_, new_G1372_, new_G1374_,
    new_G1376_, new_G1378_, new_G1380_, new_G1382_, new_G5399_, new_G5407_,
    new_G5415_, new_G5423_, new_G5431_, new_G5439_, new_G5447_, new_G5455_,
    new_G5463_, new_G5751_, new_G5759_, new_G5767_, new_G5775_, new_G5783_,
    new_G5791_, new_G5799_, new_G5807_, new_G5815_, new_G2019_, new_G2032_,
    new_G2117_, new_G2130_, new_G2266_, new_G2272_, new_G2286_, new_G2288_,
    new_G2290_, new_G2292_, new_G2294_, new_G5871_, new_G5879_, new_G5887_,
    new_G5895_, new_G5903_, new_G5911_, new_G5919_, new_G5927_, new_G5991_,
    new_G5999_, new_G6007_, new_G6015_, new_G6023_, new_G6031_, new_G6039_,
    new_G6047_, new_G2899_, new_G2914_, new_G2919_, new_G2921_, new_G2923_,
    new_G2925_, new_G2927_, new_G2929_, new_G2931_, new_G6518_, new_G3173_,
    new_G6558_, new_G6573_, new_G6581_, new_G6589_, new_G6597_, new_G6605_,
    new_G6613_, new_G6621_, new_G6629_, new_G6637_, new_G3629_, new_G3642_,
    new_G3649_, new_G3651_, new_G3653_, new_G3655_, new_G3657_, new_G3659_,
    new_G3661_, new_G3663_, new_G3762_, new_G3768_, new_G3782_, new_G3784_,
    new_G3786_, new_G3788_, new_G3790_, new_G6859_, new_G6867_, new_G6875_,
    new_G6883_, new_G6891_, new_G6899_, new_G6907_, new_G6915_, new_G6923_,
    new_G4094_, new_G4107_, new_G4444_, new_G4457_, new_G4647_, new_G4660_,
    new_G4667_, new_G4669_, new_G4671_, new_G4673_, new_G4675_, new_G4677_,
    new_G4679_, new_G4681_, new_G4683_, new_G4685_, new_G4897_, new_G5207_,
    new_G6551_, new_G763_, new_G764_, new_G4919_, new_G886_, new_G1005_,
    new_G1006_, new_G5189_, new_G1018_, new_G5237_, new_G6517_, new_G3169_,
    new_G4935_, new_G4970_, new_G5239_, new_G577_, new_G616_, new_G618_,
    new_G620_, new_G622_, new_G624_, new_G626_, new_G628_, new_G692_,
    new_G694_, new_G696_, new_G698_, new_G700_, new_G702_, new_G704_,
    new_G706_, new_G708_, new_G710_, new_G765_, new_G4903_, new_G885_,
    new_G1007_, new_G1017_, new_G5213_, new_G1363_, new_G1365_, new_G1367_,
    new_G1369_, new_G1371_, new_G1373_, new_G1375_, new_G1377_, new_G1379_,
    new_G1381_, new_G2026_, new_G2039_, new_G2046_, new_G2048_, new_G2050_,
    new_G2052_, new_G2054_, new_G2056_, new_G2058_, new_G2060_, new_G2062_,
    new_G2064_, new_G2124_, new_G2137_, new_G2144_, new_G2146_, new_G2148_,
    new_G2150_, new_G2152_, new_G2154_, new_G2156_, new_G2158_, new_G2160_,
    new_G2162_, new_G2279_, new_G2285_, new_G2287_, new_G2289_, new_G2291_,
    new_G2293_, new_G2296_, new_G2298_, new_G2300_, new_G2302_, new_G2304_,
    new_G2918_, new_G2920_, new_G2922_, new_G2924_, new_G2926_, new_G2928_,
    new_G2930_, new_G2932_, new_G3168_, new_G6557_, new_G3211_, new_G3648_,
    new_G3650_, new_G3652_, new_G3654_, new_G3656_, new_G3658_, new_G3660_,
    new_G3662_, new_G3665_, new_G3666_, new_G3775_, new_G3781_, new_G3783_,
    new_G3785_, new_G3787_, new_G3789_, new_G3792_, new_G3794_, new_G3796_,
    new_G3798_, new_G3800_, new_G4101_, new_G4114_, new_G4123_, new_G4126_,
    new_G4129_, new_G4132_, new_G4135_, new_G4138_, new_G4141_, new_G4144_,
    new_G4147_, new_G4150_, new_G4451_, new_G4464_, new_G4471_, new_G4473_,
    new_G4475_, new_G4477_, new_G4479_, new_G4481_, new_G4483_, new_G4485_,
    new_G4487_, new_G4489_, new_G4666_, new_G4668_, new_G4670_, new_G4672_,
    new_G4674_, new_G4676_, new_G4678_, new_G4680_, new_G4682_, new_G4684_,
    new_G579_, new_G629_, new_G633_, new_G637_, new_G641_, new_G645_,
    new_G711_, new_G715_, new_G719_, new_G723_, new_G727_, new_G731_,
    new_G737_, new_G745_, new_G751_, new_G757_, new_G887_, new_G1019_,
    new_G5245_, new_G1383_, new_G1387_, new_G1391_, new_G1395_, new_G1399_,
    new_G1406_, new_G1412_, new_G1418_, new_G2305_, new_G2308_, new_G2312_,
    new_G2316_, new_G2933_, new_G2938_, new_G2942_, new_G2946_, new_G2950_,
    new_G3170_, new_G3210_, new_G3667_, new_G3670_, new_G3673_, new_G3676_,
    new_G3679_, new_G3682_, new_G3686_, new_G3801_, new_G3804_, new_G3807_,
    new_G3810_, new_G3813_, new_G4525_, new_G4686_, new_G4689_, new_G4692_,
    new_G4695_, new_G4698_, new_G4701_, new_G4704_, new_G4707_, new_G4710_,
    new_G4976_, new_G5271_, new_G5274_, new_G5305_, new_G5308_, new_G5318_,
    new_G6690_, new_G6711_, new_G6714_, new_G7252_, new_G7296_, new_G7466_,
    new_G907_, new_G913_, new_G915_, new_G916_, new_G1116_, new_G2045_,
    new_G2047_, new_G2049_, new_G2051_, new_G2053_, new_G2055_, new_G2057_,
    new_G2059_, new_G2061_, new_G2063_, new_G2143_, new_G2145_, new_G2147_,
    new_G2149_, new_G2151_, new_G2153_, new_G2155_, new_G2157_, new_G2159_,
    new_G2161_, new_G2295_, new_G2297_, new_G2299_, new_G2301_, new_G2303_,
    new_G3212_, new_G3791_, new_G3793_, new_G3795_, new_G3797_, new_G3799_,
    new_G4122_, new_G4125_, new_G4128_, new_G4131_, new_G4134_, new_G4137_,
    new_G4140_, new_G4143_, new_G4146_, new_G4149_, new_G4470_, new_G4472_,
    new_G4474_, new_G4476_, new_G4478_, new_G4480_, new_G4482_, new_G4484_,
    new_G4486_, new_G4488_, new_G4962_, new_G5003_, new_G5234_, new_G5242_,
    new_G5250_, new_G5284_, new_G802_, new_G821_, new_G845_, new_G868_,
    new_G877_, new_G902_, new_G908_, new_G914_, new_G917_, new_G953_,
    new_G1023_, new_G1035_, new_G1050_, new_G1068_, new_G1086_, new_G1102_,
    new_G1108_, new_G1117_, new_G5322_, new_G1553_, new_G1567_, new_G1584_,
    new_G1590_, new_G1606_, new_G1624_, new_G1647_, new_G1669_, new_G1677_,
    new_G1802_, new_G1816_, new_G1834_, new_G1841_, new_G1866_, new_G1880_,
    new_G1897_, new_G1914_, new_G1929_, new_G2065_, new_G2069_, new_G2073_,
    new_G2077_, new_G2081_, new_G2085_, new_G2091_, new_G2099_, new_G2105_,
    new_G2111_, new_G2163_, new_G2167_, new_G2171_, new_G2175_, new_G2179_,
    new_G2186_, new_G2192_, new_G2198_, new_G2320_, new_G2323_, new_G2329_,
    new_G2335_, new_G2962_, new_G2970_, new_G2977_, new_G2979_, new_G2989_,
    new_G2998_, new_G3006_, new_G3013_, new_G3015_, new_G3183_, new_G3192_,
    new_G3200_, new_G3207_, new_G3209_, new_G3216_, new_G3222_, new_G6694_,
    new_G3695_, new_G3816_, new_G3821_, new_G3828_, new_G3833_, new_G3838_,
    new_G4151_, new_G4154_, new_G4157_, new_G4160_, new_G4163_, new_G4166_,
    new_G4169_, new_G4172_, new_G4175_, new_G7256_, new_G7300_, new_G4490_,
    new_G4493_, new_G4496_, new_G4499_, new_G4502_, new_G4505_, new_G4508_,
    new_G4511_, new_G7470_, new_G4884_, new_G4892_, new_G4900_, new_G4908_,
    new_G4924_, new_G4952_, new_G4983_, new_G4993_, new_G5011_, new_G5194_,
    new_G5202_, new_G5210_, new_G5218_, new_G5226_, new_G5247_, new_G5255_,
    new_G5258_, new_G5263_, new_G5266_, new_G5277_, new_G5278_, new_G5281_,
    new_G5289_, new_G5292_, new_G5297_, new_G5300_, new_G5311_, new_G5312_,
    new_G5315_, new_G5323_, new_G5326_, new_G5331_, new_G5334_, new_G5339_,
    new_G5342_, new_G5349_, new_G5352_, new_G5396_, new_G5404_, new_G5412_,
    new_G5420_, new_G5428_, new_G5436_, new_G5444_, new_G5452_, new_G5460_,
    new_G5465_, new_G5581_, new_G5748_, new_G5756_, new_G5764_, new_G5772_,
    new_G5780_, new_G5788_, new_G5796_, new_G5804_, new_G5812_, new_G5849_,
    new_G5929_, new_G6049_, new_G6367_, new_G6370_, new_G6375_, new_G6378_,
    new_G6383_, new_G6386_, new_G6391_, new_G6394_, new_G6399_, new_G6402_,
    new_G6407_, new_G6410_, new_G6415_, new_G6418_, new_G6423_, new_G6426_,
    new_G6431_, new_G6434_, new_G6442_, new_G6450_, new_G6458_, new_G6466_,
    new_G6498_, new_G6519_, new_G6522_, new_G6527_, new_G6530_, new_G6535_,
    new_G6538_, new_G6543_, new_G6546_, new_G6559_, new_G6562_, new_G6687_,
    new_G6695_, new_G6698_, new_G6703_, new_G6706_, new_G6717_, new_G6718_,
    new_G6724_, new_G6768_, new_G7208_, new_G7221_, new_G7229_, new_G7232_,
    new_G7239_, new_G7242_, new_G7249_, new_G7257_, new_G7260_, new_G7268_,
    new_G7293_, new_G7301_, new_G7304_, new_G7309_, new_G7312_, new_G7317_,
    new_G7320_, new_G7327_, new_G7330_, new_G7396_, new_G7404_, new_G7412_,
    new_G7425_, new_G7463_, new_G7471_, new_G7474_, new_G7479_, new_G7482_,
    new_G7487_, new_G7490_, new_G7497_, new_G7500_, new_G7507_, new_G7510_,
    new_G7554_, new_G1152_, new_G5238_, new_G1156_, new_G5246_, new_G5254_,
    new_G5288_, new_G3223_, new_G4942_, new_G4966_, new_G5007_, new_G5279_,
    new_G5280_, new_G5313_, new_G5314_, new_G6719_, new_G6720_, new_G790_,
    new_G4888_, new_G803_, new_G4896_, new_G825_, new_G4904_, new_G851_,
    new_G4912_, new_G893_, new_G4928_, new_G906_, new_G912_, new_G1024_,
    new_G5198_, new_G1036_, new_G5206_, new_G1053_, new_G5214_, new_G1072_,
    new_G5222_, new_G1091_, new_G5230_, new_G1112_, new_G1121_, new_G1153_,
    new_G1157_, new_G5253_, new_G1216_, new_G5261_, new_G5262_, new_G5269_,
    new_G5270_, new_G5287_, new_G1239_, new_G5295_, new_G5296_, new_G5303_,
    new_G5304_, new_G5321_, new_G1262_, new_G5329_, new_G5330_, new_G5337_,
    new_G5338_, new_G1544_, new_G5400_, new_G1554_, new_G5408_, new_G1571_,
    new_G5416_, new_G1596_, new_G5424_, new_G1607_, new_G5432_, new_G1628_,
    new_G5440_, new_G1653_, new_G5448_, new_G1685_, new_G5456_, new_G1693_,
    new_G5464_, new_G1793_, new_G5752_, new_G1803_, new_G5760_, new_G1820_,
    new_G5768_, new_G1848_, new_G5776_, new_G1857_, new_G5784_, new_G1867_,
    new_G5792_, new_G1883_, new_G5800_, new_G1901_, new_G5808_, new_G1919_,
    new_G5816_, new_G5855_, new_G2351_, new_G2366_, new_G2384_, new_G2391_,
    new_G2417_, new_G2431_, new_G2448_, new_G2465_, new_G5935_, new_G2597_,
    new_G2612_, new_G2629_, new_G2635_, new_G2652_, new_G2670_, new_G2693_,
    new_G2715_, new_G6055_, new_G6373_, new_G6374_, new_G6381_, new_G6382_,
    new_G6389_, new_G6390_, new_G6397_, new_G6398_, new_G6405_, new_G6406_,
    new_G6413_, new_G6414_, new_G6421_, new_G6422_, new_G6429_, new_G6430_,
    new_G6437_, new_G6438_, new_G6446_, new_G3059_, new_G6454_, new_G3068_,
    new_G6462_, new_G3076_, new_G3079_, new_G6470_, new_G3090_, new_G3099_,
    new_G3107_, new_G3114_, new_G3116_, new_G6502_, new_G6525_, new_G6526_,
    new_G6533_, new_G6534_, new_G6541_, new_G6542_, new_G6549_, new_G6550_,
    new_G6565_, new_G6566_, new_G3220_, new_G3292_, new_G3308_, new_G3327_,
    new_G3335_, new_G3362_, new_G3376_, new_G3393_, new_G3410_, new_G3425_,
    new_G6693_, new_G3503_, new_G6701_, new_G6702_, new_G6709_, new_G6710_,
    new_G6728_, new_G6772_, new_G3853_, new_G3868_, new_G3885_, new_G3891_,
    new_G3908_, new_G3926_, new_G3949_, new_G3971_, new_G3979_, new_G7212_,
    new_G7227_, new_G7255_, new_G4202_, new_G7263_, new_G7264_, new_G7272_,
    new_G7299_, new_G4225_, new_G7307_, new_G7308_, new_G7315_, new_G7316_,
    new_G4297_, new_G4305_, new_G4312_, new_G4314_, new_G4324_, new_G7400_,
    new_G4333_, new_G7408_, new_G4341_, new_G7416_, new_G4348_, new_G4349_,
    new_G7431_, new_G4389_, new_G7469_, new_G4530_, new_G7477_, new_G7478_,
    new_G7485_, new_G7486_, new_G7513_, new_G7514_, new_G7558_, new_G4932_,
    new_G4956_, new_G4973_, new_G4987_, new_G4997_, new_G5017_, new_G5099_,
    new_G5345_, new_G5346_, new_G5355_, new_G5356_, new_G5372_, new_G5380_,
    new_G5471_, new_G5523_, new_G5587_, new_G5669_, new_G5857_, new_G5868_,
    new_G5876_, new_G5884_, new_G5892_, new_G5900_, new_G5908_, new_G5916_,
    new_G5924_, new_G5969_, new_G5988_, new_G5996_, new_G6004_, new_G6012_,
    new_G6020_, new_G6028_, new_G6036_, new_G6044_, new_G6057_, new_G6439_,
    new_G6447_, new_G6455_, new_G6463_, new_G6471_, new_G6474_, new_G6479_,
    new_G6482_, new_G6487_, new_G6490_, new_G6495_, new_G6503_, new_G6506_,
    new_G6570_, new_G6578_, new_G6586_, new_G6594_, new_G6602_, new_G6610_,
    new_G6618_, new_G6626_, new_G6634_, new_G6671_, new_G6721_, new_G6729_,
    new_G6732_, new_G6737_, new_G6740_, new_G6745_, new_G6748_, new_G6755_,
    new_G6758_, new_G6765_, new_G6773_, new_G6776_, new_G6781_, new_G6784_,
    new_G6789_, new_G6792_, new_G6799_, new_G6802_, new_G6832_, new_G6856_,
    new_G6864_, new_G6872_, new_G6880_, new_G6888_, new_G6896_, new_G6904_,
    new_G6912_, new_G6920_, new_G6925_, new_G7041_, new_G7205_, new_G7213_,
    new_G7216_, new_G7224_, new_G7235_, new_G7236_, new_G7245_, new_G7246_,
    new_G7265_, new_G7273_, new_G7276_, new_G7283_, new_G7286_, new_G7323_,
    new_G7324_, new_G7333_, new_G7334_, new_G7361_, new_G7364_, new_G7369_,
    new_G7372_, new_G7377_, new_G7380_, new_G7385_, new_G7388_, new_G7393_,
    new_G7401_, new_G7409_, new_G7417_, new_G7420_, new_G7428_, new_G7493_,
    new_G7494_, new_G7503_, new_G7504_, new_G7515_, new_G7518_, new_G7523_,
    new_G7526_, new_G7531_, new_G7534_, new_G7541_, new_G7544_, new_G7551_,
    new_G7559_, new_G7562_, new_G7567_, new_G7570_, new_G7575_, new_G7578_,
    new_G7585_, new_G7588_, new_G1176_, new_G957_, new_G791_, new_G804_,
    new_G826_, new_G852_, new_G894_, new_G1025_, new_G1037_, new_G1054_,
    new_G1073_, new_G1092_, new_G1154_, new_G1158_, new_G1215_, new_G1224_,
    new_G1225_, new_G1233_, new_G1234_, new_G1238_, new_G1247_, new_G1248_,
    new_G1256_, new_G1257_, new_G1261_, new_G1270_, new_G1271_, new_G1279_,
    new_G1280_, new_G1545_, new_G1555_, new_G1572_, new_G1597_, new_G1608_,
    new_G1629_, new_G1654_, new_G1686_, new_G1694_, new_G1794_, new_G1804_,
    new_G1821_, new_G1849_, new_G1858_, new_G1868_, new_G1884_, new_G1902_,
    new_G1920_, new_G2954_, new_G2955_, new_G2963_, new_G2964_, new_G2971_,
    new_G2972_, new_G2980_, new_G2981_, new_G2990_, new_G2991_, new_G2999_,
    new_G3000_, new_G3007_, new_G3008_, new_G3016_, new_G3017_, new_G3019_,
    new_G3020_, new_G3174_, new_G3175_, new_G3184_, new_G3185_, new_G3193_,
    new_G3194_, new_G3201_, new_G3202_, new_G3213_, new_G3214_, new_G3227_,
    new_G3502_, new_G3511_, new_G3512_, new_G3520_, new_G3521_, new_G4201_,
    new_G4210_, new_G4211_, new_G4224_, new_G4233_, new_G4234_, new_G4242_,
    new_G4243_, new_G4529_, new_G4538_, new_G4539_, new_G4547_, new_G4548_,
    new_G4552_, new_G4553_, new_G4946_, new_G5347_, new_G5348_, new_G5357_,
    new_G5358_, new_G7237_, new_G7238_, new_G7247_, new_G7248_, new_G7325_,
    new_G7326_, new_G7335_, new_G7336_, new_G7495_, new_G7496_, new_G7505_,
    new_G7506_, new_G3244_, new_G792_, new_G805_, new_G827_, new_G853_,
    new_G895_, new_G1026_, new_G1038_, new_G1055_, new_G1074_, new_G1093_,
    new_G1155_, new_G1217_, new_G1226_, new_G1235_, new_G1240_, new_G1249_,
    new_G1258_, new_G1263_, new_G1272_, new_G1281_, new_G5376_, new_G5384_,
    new_G1546_, new_G1556_, new_G1573_, new_G1598_, new_G1609_, new_G1630_,
    new_G1655_, new_G1687_, new_G1695_, new_G1795_, new_G1805_, new_G1822_,
    new_G1850_, new_G1859_, new_G1869_, new_G1885_, new_G1903_, new_G1921_,
    new_G5863_, new_G2341_, new_G5872_, new_G2352_, new_G5880_, new_G2370_,
    new_G5888_, new_G2398_, new_G5896_, new_G2407_, new_G5904_, new_G2418_,
    new_G5912_, new_G2434_, new_G5920_, new_G2452_, new_G5928_, new_G2481_,
    new_G5975_, new_G2587_, new_G5992_, new_G2598_, new_G6000_, new_G2616_,
    new_G6008_, new_G2641_, new_G6016_, new_G2653_, new_G6024_, new_G2674_,
    new_G6032_, new_G2699_, new_G6040_, new_G2724_, new_G2732_, new_G6048_,
    new_G2956_, new_G2965_, new_G2973_, new_G2982_, new_G2992_, new_G3001_,
    new_G3009_, new_G3018_, new_G3021_, new_G6445_, new_G3051_, new_G6453_,
    new_G3061_, new_G6461_, new_G3070_, new_G6469_, new_G3081_, new_G6477_,
    new_G6478_, new_G6485_, new_G6486_, new_G6493_, new_G6494_, new_G6501_,
    new_G3118_, new_G6509_, new_G6510_, new_G3176_, new_G3186_, new_G3195_,
    new_G3203_, new_G3215_, new_G3281_, new_G6574_, new_G3293_, new_G6582_,
    new_G3312_, new_G6590_, new_G3342_, new_G6598_, new_G3351_, new_G6606_,
    new_G3363_, new_G6614_, new_G3379_, new_G6622_, new_G3397_, new_G6630_,
    new_G3415_, new_G6638_, new_G6677_, new_G3504_, new_G3513_, new_G3522_,
    new_G6727_, new_G3526_, new_G6735_, new_G6736_, new_G6743_, new_G6744_,
    new_G6771_, new_G3549_, new_G6779_, new_G6780_, new_G6787_, new_G6788_,
    new_G6836_, new_G3843_, new_G6860_, new_G3854_, new_G6868_, new_G3872_,
    new_G6876_, new_G3897_, new_G6884_, new_G3909_, new_G6892_, new_G3930_,
    new_G6900_, new_G3955_, new_G6908_, new_G3987_, new_G6916_, new_G3995_,
    new_G6924_, new_G7211_, new_G4179_, new_G7219_, new_G7220_, new_G4196_,
    new_G7228_, new_G4203_, new_G4212_, new_G7271_, new_G4220_, new_G4226_,
    new_G4235_, new_G4244_, new_G7367_, new_G7368_, new_G7375_, new_G7376_,
    new_G7383_, new_G7384_, new_G7391_, new_G7392_, new_G7399_, new_G4326_,
    new_G7407_, new_G4335_, new_G7415_, new_G4343_, new_G7423_, new_G7424_,
    new_G4353_, new_G7432_, new_G4531_, new_G4540_, new_G4549_, new_G4554_,
    new_G7521_, new_G7522_, new_G7529_, new_G7530_, new_G7557_, new_G4576_,
    new_G7565_, new_G7566_, new_G7573_, new_G7574_, new_G4936_, new_G4937_,
    new_G4977_, new_G4978_, new_G5105_, new_G5359_, new_G5362_, new_G5529_,
    new_G5675_, new_G5932_, new_G5977_, new_G6052_, new_G6063_, new_G6115_,
    new_G6173_, new_G6679_, new_G6751_, new_G6752_, new_G6761_, new_G6762_,
    new_G6795_, new_G6796_, new_G6805_, new_G6806_, new_G6931_, new_G6983_,
    new_G7047_, new_G7129_, new_G7279_, new_G7280_, new_G7289_, new_G7290_,
    new_G7337_, new_G7340_, new_G7353_, new_G7356_, new_G7537_, new_G7538_,
    new_G7547_, new_G7548_, new_G7581_, new_G7582_, new_G7591_, new_G7592_,
    new_G7595_, new_G7598_, new_G2342_, new_G2353_, new_G2371_, new_G2399_,
    new_G2408_, new_G2419_, new_G2435_, new_G2453_, new_G2588_, new_G2599_,
    new_G2617_, new_G2642_, new_G2654_, new_G2675_, new_G2700_, new_G2733_,
    new_G3050_, new_G3060_, new_G3069_, new_G3080_, new_G3091_, new_G3092_,
    new_G3100_, new_G3101_, new_G3108_, new_G3109_, new_G3117_, new_G3120_,
    new_G3121_, new_G3282_, new_G3294_, new_G3313_, new_G3343_, new_G3352_,
    new_G3364_, new_G3380_, new_G3398_, new_G3416_, new_G3525_, new_G3534_,
    new_G3535_, new_G3543_, new_G3544_, new_G3548_, new_G3557_, new_G3558_,
    new_G3566_, new_G3567_, new_G3844_, new_G3855_, new_G3873_, new_G3898_,
    new_G3910_, new_G3931_, new_G3956_, new_G3988_, new_G3996_, new_G4178_,
    new_G4187_, new_G4188_, new_G4197_, new_G4219_, new_G4289_, new_G4290_,
    new_G4298_, new_G4299_, new_G4306_, new_G4307_, new_G4315_, new_G4316_,
    new_G4325_, new_G4334_, new_G4342_, new_G4350_, new_G4351_, new_G4354_,
    new_G4561_, new_G4562_, new_G4570_, new_G4571_, new_G4575_, new_G4584_,
    new_G4585_, new_G4593_, new_G4594_, new_G4938_, new_G4979_, new_G6753_,
    new_G6754_, new_G6763_, new_G6764_, new_G6797_, new_G6798_, new_G6807_,
    new_G6808_, new_G7281_, new_G7282_, new_G7291_, new_G7292_, new_G7539_,
    new_G7540_, new_G7549_, new_G7550_, new_G7583_, new_G7584_, new_G7593_,
    new_G7594_, new_G1856_, new_G920_, new_G925_, new_G926_, new_G927_,
    new_G928_, new_G937_, new_G938_, new_G939_, new_G940_, new_G941_,
    new_G942_, new_G943_, new_G944_, new_G945_, new_G946_, new_G947_,
    new_G948_, new_G949_, new_G956_, new_G1122_, new_G1125_, new_G1126_,
    new_G1127_, new_G1128_, new_G1132_, new_G1133_, new_G1134_, new_G1137_,
    new_G1138_, new_G1141_, new_G1221_, new_G1230_, new_G1244_, new_G1253_,
    new_G1267_, new_G1276_, new_G1284_, new_G1288_, new_G1292_, new_G1296_,
    new_G1300_, new_G1304_, new_G1702_, new_G1705_, new_G1706_, new_G1707_,
    new_G1709_, new_G1710_, new_G1711_, new_G1712_, new_G1713_, new_G1714_,
    new_G1718_, new_G1722_, new_G1723_, new_G1724_, new_G1725_, new_G1733_,
    new_G1734_, new_G1735_, new_G1736_, new_G1737_, new_G1738_, new_G1739_,
    new_G1740_, new_G1741_, new_G1742_, new_G1743_, new_G1744_, new_G1745_,
    new_G1749_, new_G1750_, new_G1935_, new_G1938_, new_G1939_, new_G1940_,
    new_G1942_, new_G1943_, new_G1944_, new_G1945_, new_G1946_, new_G1947_,
    new_G1948_, new_G1949_, new_G1950_, new_G1953_, new_G1954_, new_G1955_,
    new_G1956_, new_G1960_, new_G1961_, new_G1962_, new_G1965_, new_G1966_,
    new_G1969_, new_G2343_, new_G2354_, new_G2372_, new_G2400_, new_G2409_,
    new_G2420_, new_G2436_, new_G2454_, new_G2470_, new_G5936_, new_G5983_,
    new_G2589_, new_G2600_, new_G2618_, new_G2643_, new_G2655_, new_G2676_,
    new_G2701_, new_G2734_, new_G2740_, new_G6056_, new_G3022_, new_G3025_,
    new_G3026_, new_G3027_, new_G3029_, new_G3030_, new_G3031_, new_G3032_,
    new_G3033_, new_G3052_, new_G3062_, new_G3071_, new_G3082_, new_G3093_,
    new_G3102_, new_G3110_, new_G3119_, new_G3122_, new_G3228_, new_G3231_,
    new_G3232_, new_G3233_, new_G3234_, new_G3283_, new_G3295_, new_G3314_,
    new_G3344_, new_G3353_, new_G3365_, new_G3381_, new_G3399_, new_G3417_,
    new_G6685_, new_G3508_, new_G3517_, new_G3527_, new_G3536_, new_G3545_,
    new_G3550_, new_G3559_, new_G3568_, new_G3571_, new_G3575_, new_G3845_,
    new_G3856_, new_G3874_, new_G3899_, new_G3911_, new_G3932_, new_G3957_,
    new_G3989_, new_G3997_, new_G4180_, new_G4189_, new_G4198_, new_G4207_,
    new_G4216_, new_G4221_, new_G4230_, new_G4239_, new_G4263_, new_G4267_,
    new_G4291_, new_G4300_, new_G4308_, new_G4317_, new_G4327_, new_G4336_,
    new_G4344_, new_G4352_, new_G4355_, new_G4535_, new_G4544_, new_G4558_,
    new_G4563_, new_G4572_, new_G4577_, new_G4586_, new_G4595_, new_G4598_,
    new_G4602_, new_G4716_, new_G4724_, new_G4732_, new_G4740_, new_G4748_,
    new_G4756_, new_G4764_, new_G4772_, new_G4780_, new_G4788_, new_G4939_,
    new_G4980_, new_G5044_, new_G5054_, new_G5064_, new_G5074_, new_G5084_,
    new_G5094_, new_G5132_, new_G5142_, new_G5152_, new_G5162_, new_G5365_,
    new_G5366_, new_G5488_, new_G5498_, new_G5508_, new_G5518_, new_G5546_,
    new_G5556_, new_G5566_, new_G5576_, new_G5614_, new_G5624_, new_G5634_,
    new_G5644_, new_G5654_, new_G5664_, new_G5702_, new_G5712_, new_G5722_,
    new_G5732_, new_G5820_, new_G5828_, new_G5836_, new_G5844_, new_G5852_,
    new_G5860_, new_G6121_, new_G6179_, new_G6261_, new_G7359_, new_G7360_,
    new_G7343_, new_G7344_, new_G6809_, new_G6812_, new_G6819_, new_G6822_,
    new_G6989_, new_G7135_, new_G7345_, new_G7348_, new_G7601_, new_G7602_,
    new_G7603_, new_G7606_, new_G7611_, new_G7614_, new_G929_, new_G950_,
    new_G1129_, new_G1708_, new_G1715_, new_G1726_, new_G1746_, new_G1941_,
    new_G1957_, new_G2471_, new_G2741_, new_G3028_, new_G3034_, new_G3235_,
    new_G5014_, new_G5034_, new_G5102_, new_G5122_, new_G5367_, new_G5368_,
    new_G5478_, new_G5536_, new_G5584_, new_G5604_, new_G5672_, new_G5692_,
    new_G5817_, new_G5825_, new_G5833_, new_G5841_, new_G6340_, new_G6341_,
    new_G6350_, new_G6351_, new_G7436_, new_G7437_, new_G4720_, new_G4728_,
    new_G4736_, new_G4744_, new_G4752_, new_G4760_, new_G4768_, new_G4776_,
    new_G4784_, new_G4792_, new_G3350_, new_G2406_, new_G924_, new_G5088_,
    new_G5098_, new_G997_, new_G1146_, new_G1287_, new_G1291_, new_G1295_,
    new_G1299_, new_G1303_, new_G1307_, new_G1309_, new_G1312_, new_G1315_,
    new_G1318_, new_G1321_, new_G1324_, new_G1721_, new_G5522_, new_G5580_,
    new_G5658_, new_G5668_, new_G1788_, new_G1974_, new_G5824_, new_G5832_,
    new_G5840_, new_G5848_, new_G1999_, new_G5856_, new_G2003_, new_G5864_,
    new_G2472_, new_G2487_, new_G2492_, new_G2493_, new_G2494_, new_G2500_,
    new_G2501_, new_G2502_, new_G2503_, new_G2504_, new_G2505_, new_G2506_,
    new_G2507_, new_G2511_, new_G2512_, new_G2513_, new_G2514_, new_G2518_,
    new_G2519_, new_G2520_, new_G2523_, new_G2524_, new_G2527_, new_G2742_,
    new_G2749_, new_G2754_, new_G2755_, new_G2756_, new_G2762_, new_G2763_,
    new_G2764_, new_G2765_, new_G2766_, new_G2767_, new_G2776_, new_G2777_,
    new_G2778_, new_G2779_, new_G2788_, new_G2789_, new_G2790_, new_G2792_,
    new_G2793_, new_G2794_, new_G2795_, new_G2796_, new_G2798_, new_G2799_,
    new_G2800_, new_G2804_, new_G3035_, new_G3045_, new_G3123_, new_G3128_,
    new_G3129_, new_G3130_, new_G3136_, new_G3139_, new_G3140_, new_G3141_,
    new_G3142_, new_G3249_, new_G3431_, new_G3434_, new_G3435_, new_G3436_,
    new_G3438_, new_G3439_, new_G3440_, new_G3441_, new_G3442_, new_G3443_,
    new_G3444_, new_G3445_, new_G3446_, new_G3449_, new_G3450_, new_G3451_,
    new_G3452_, new_G3456_, new_G3457_, new_G3458_, new_G3460_, new_G3461_,
    new_G3463_, new_G3531_, new_G3540_, new_G3554_, new_G3563_, new_G3574_,
    new_G3578_, new_G3579_, new_G3583_, new_G3587_, new_G3591_, new_G3596_,
    new_G3599_, new_G4004_, new_G4007_, new_G4008_, new_G4009_, new_G4011_,
    new_G4012_, new_G4013_, new_G4014_, new_G4015_, new_G4016_, new_G4020_,
    new_G4024_, new_G4025_, new_G4026_, new_G4027_, new_G4035_, new_G4036_,
    new_G4037_, new_G4038_, new_G4039_, new_G4040_, new_G4041_, new_G4042_,
    new_G4043_, new_G4044_, new_G4045_, new_G4046_, new_G4047_, new_G4051_,
    new_G4052_, new_G4184_, new_G4193_, new_G4247_, new_G4251_, new_G4255_,
    new_G4259_, new_G4266_, new_G4270_, new_G4284_, new_G4287_, new_G4356_,
    new_G4361_, new_G4362_, new_G4363_, new_G4369_, new_G4372_, new_G4373_,
    new_G4374_, new_G4375_, new_G4567_, new_G4581_, new_G4590_, new_G4601_,
    new_G4605_, new_G4606_, new_G4610_, new_G4614_, new_G4618_, new_G4623_,
    new_G4626_, new_G4796_, new_G4804_, new_G4812_, new_G4820_, new_G4828_,
    new_G4844_, new_G4852_, new_G4860_, new_G4868_, new_G4945_, new_G4948_,
    new_G4986_, new_G4989_, new_G5048_, new_G5058_, new_G5068_, new_G5078_,
    new_G5166_, new_G5136_, new_G5146_, new_G5156_, new_G5388_, new_G5492_,
    new_G5502_, new_G5512_, new_G5550_, new_G5560_, new_G5570_, new_G5618_,
    new_G5628_, new_G5638_, new_G5648_, new_G5736_, new_G5706_, new_G5716_,
    new_G5726_, new_G5940_, new_G5948_, new_G5956_, new_G5964_, new_G5972_,
    new_G5980_, new_G6080_, new_G6090_, new_G6100_, new_G6110_, new_G6138_,
    new_G6148_, new_G6158_, new_G6168_, new_G6216_, new_G6226_, new_G6236_,
    new_G6246_, new_G6256_, new_G6267_, new_G6304_, new_G6314_, new_G6324_,
    new_G6342_, new_G6352_, new_G7351_, new_G7352_, new_G6642_, new_G6650_,
    new_G6658_, new_G6666_, new_G6674_, new_G6682_, new_G6815_, new_G6816_,
    new_G6825_, new_G6826_, new_G6948_, new_G6958_, new_G6968_, new_G6978_,
    new_G7006_, new_G7016_, new_G7026_, new_G7036_, new_G7074_, new_G7084_,
    new_G7094_, new_G7104_, new_G7114_, new_G7124_, new_G7162_, new_G7172_,
    new_G7182_, new_G7192_, new_G7438_, new_G7617_, new_G7618_, new_G7609_,
    new_G7610_, new_G1151_, new_G1002_, new_G933_, new_G1308_, new_G1311_,
    new_G1314_, new_G1317_, new_G1320_, new_G1323_, new_G1730_, new_G1789_,
    new_G1981_, new_G5823_, new_G1986_, new_G5831_, new_G1989_, new_G5839_,
    new_G1993_, new_G5847_, new_G1996_, new_G2000_, new_G2004_, new_G2495_,
    new_G2515_, new_G2757_, new_G2768_, new_G2780_, new_G2801_, new_G3046_,
    new_G3131_, new_G3143_, new_G3238_, new_G3258_, new_G3437_, new_G3453_,
    new_G3595_, new_G3598_, new_G4010_, new_G4017_, new_G4028_, new_G4048_,
    new_G4283_, new_G4286_, new_G4364_, new_G4376_, new_G4622_, new_G4625_,
    new_G4947_, new_G4988_, new_G5018_, new_G5019_, new_G5024_, new_G5038_,
    new_G5106_, new_G5107_, new_G5112_, new_G5126_, new_G5468_, new_G5482_,
    new_G5526_, new_G5540_, new_G5588_, new_G5589_, new_G5594_, new_G5608_,
    new_G5676_, new_G5677_, new_G5682_, new_G5696_, new_G5937_, new_G5945_,
    new_G5953_, new_G5961_, new_G6070_, new_G6128_, new_G6264_, new_G6284_,
    new_G6360_, new_G6361_, new_G6639_, new_G6647_, new_G6655_, new_G6663_,
    new_G6817_, new_G6818_, new_G6827_, new_G6828_, new_G6938_, new_G6996_,
    new_G7044_, new_G7064_, new_G7132_, new_G7152_, new_G7446_, new_G7447_,
    new_G7456_, new_G7457_, new_G241_, new_G265_, new_G2005_, new_G4800_,
    new_G4808_, new_G4816_, new_G4824_, new_G4832_, new_G4848_, new_G4856_,
    new_G4864_, new_G4872_, new_G1310_, new_G1313_, new_G1316_, new_G1319_,
    new_G1322_, new_G1325_, new_G5392_, new_G1790_, new_G1982_, new_G1985_,
    new_G1988_, new_G1992_, new_G1995_, new_G2001_, new_G2491_, new_G2508_,
    new_G2522_, new_G2526_, new_G2529_, new_G2531_, new_G5944_, new_G5952_,
    new_G5960_, new_G5968_, new_G2555_, new_G5976_, new_G2559_, new_G5984_,
    new_G2753_, new_G2771_, new_G2791_, new_G2797_, new_G2807_, new_G6114_,
    new_G6172_, new_G6250_, new_G6260_, new_G6346_, new_G6356_, new_G3127_,
    new_G3156_, new_G3259_, new_G3466_, new_G6646_, new_G6654_, new_G6662_,
    new_G6670_, new_G3483_, new_G6678_, new_G3487_, new_G6686_, new_G3582_,
    new_G3586_, new_G3590_, new_G3594_, new_G3597_, new_G3600_, new_G3602_,
    new_G3605_, new_G3608_, new_G3611_, new_G4023_, new_G6982_, new_G7040_,
    new_G7118_, new_G7128_, new_G4089_, new_G4250_, new_G4254_, new_G4258_,
    new_G4262_, new_G4272_, new_G4275_, new_G4278_, new_G4281_, new_G4285_,
    new_G4288_, new_G4360_, new_G4380_, new_G4386_, new_G7442_, new_G4609_,
    new_G4613_, new_G4617_, new_G4621_, new_G4624_, new_G4627_, new_G4629_,
    new_G4632_, new_G4635_, new_G4638_, new_G4836_, new_G4949_, new_G4990_,
    new_G5020_, new_G5108_, new_G5590_, new_G5678_, new_G6084_, new_G6094_,
    new_G6104_, new_G6142_, new_G6152_, new_G6162_, new_G6206_, new_G6220_,
    new_G6230_, new_G6240_, new_G6328_, new_G6294_, new_G6308_, new_G6318_,
    new_G6362_, new_G6840_, new_G6848_, new_G6952_, new_G6962_, new_G6972_,
    new_G7010_, new_G7020_, new_G7030_, new_G7078_, new_G7088_, new_G7098_,
    new_G7108_, new_G7196_, new_G7166_, new_G7176_, new_G7186_, new_G7448_,
    new_G7458_, new_G254_, new_G260_, new_G1987_, new_G1994_, new_G2002_,
    new_G962_, new_G1751_, new_G1990_, new_G1997_, new_G2499_, new_G2536_,
    new_G5943_, new_G2542_, new_G5951_, new_G2545_, new_G5959_, new_G2549_,
    new_G5967_, new_G2552_, new_G2556_, new_G2560_, new_G2761_, new_G2784_,
    new_G2853_, new_G3135_, new_G3146_, new_G3163_, new_G3467_, new_G6645_,
    new_G3470_, new_G6653_, new_G3473_, new_G6661_, new_G3477_, new_G6669_,
    new_G3480_, new_G3484_, new_G3488_, new_G3601_, new_G3604_, new_G3607_,
    new_G3610_, new_G4032_, new_G4090_, new_G4271_, new_G4274_, new_G4277_,
    new_G4280_, new_G4368_, new_G4379_, new_G4387_, new_G4628_, new_G4631_,
    new_G4634_, new_G4637_, new_G4841_, new_G4849_, new_G4857_, new_G4865_,
    new_G5021_, new_G5028_, new_G5109_, new_G5116_, new_G5369_, new_G5377_,
    new_G5385_, new_G5472_, new_G5473_, new_G5530_, new_G5531_, new_G5591_,
    new_G5598_, new_G5679_, new_G5686_, new_G6060_, new_G6074_, new_G6118_,
    new_G6132_, new_G6176_, new_G6186_, new_G6196_, new_G6268_, new_G6269_,
    new_G6274_, new_G6288_, new_G6337_, new_G6829_, new_G6928_, new_G6942_,
    new_G6986_, new_G7000_, new_G7048_, new_G7049_, new_G7054_, new_G7068_,
    new_G7136_, new_G7137_, new_G7142_, new_G7156_, new_G7433_, new_G242_,
    new_G3151_, new_G257_, new_G263_, new_G266_, new_G1991_, new_G1998_,
    new_G3489_, new_G371_, new_G4840_, new_G2561_, new_G2532_, new_G2537_,
    new_G2541_, new_G2544_, new_G2548_, new_G2551_, new_G2557_, new_G2563_,
    new_G2577_, new_G2775_, new_G2806_, new_G2808_, new_G2852_, new_G2854_,
    new_G6366_, new_G4381_, new_G3164_, new_G3241_, new_G3468_, new_G3469_,
    new_G3472_, new_G3476_, new_G3479_, new_G3485_, new_G3603_, new_G3606_,
    new_G3609_, new_G3612_, new_G6844_, new_G6852_, new_G4091_, new_G4273_,
    new_G4276_, new_G4279_, new_G4282_, new_G4382_, new_G4388_, new_G7452_,
    new_G7462_, new_G4630_, new_G4633_, new_G4636_, new_G4639_, new_G4955_,
    new_G4958_, new_G4996_, new_G4999_, new_G5474_, new_G5532_, new_G6210_,
    new_G6270_, new_G6298_, new_G7050_, new_G7138_, new_G3471_, new_G3478_,
    new_G3486_, new_G372_, new_G2543_, new_G2550_, new_G2558_, new_G4847_,
    new_G387_, new_G4855_, new_G390_, new_G4863_, new_G393_, new_G4871_,
    new_G396_, new_G965_, new_G5375_, new_G1327_, new_G5383_, new_G1330_,
    new_G5391_, new_G1333_, new_G1754_, new_G2546_, new_G2553_, new_G2564_,
    new_G2809_, new_G2813_, new_G6345_, new_G2860_, new_G3474_, new_G3481_,
    new_G6835_, new_G3614_, new_G4053_, new_G7441_, new_G4516_, new_G4957_,
    new_G4998_, new_G5027_, new_G5030_, new_G5115_, new_G5118_, new_G5475_,
    new_G5533_, new_G5597_, new_G5600_, new_G5685_, new_G5688_, new_G6064_,
    new_G6065_, new_G6122_, new_G6123_, new_G6180_, new_G6181_, new_G6190_,
    new_G6200_, new_G6271_, new_G6278_, new_G6347_, new_G6357_, new_G6837_,
    new_G6845_, new_G6932_, new_G6933_, new_G6990_, new_G6991_, new_G7051_,
    new_G7058_, new_G7139_, new_G7146_, new_G7443_, new_G7453_, new_G243_,
    new_G244_, new_G245_, new_G255_, new_G256_, new_G261_, new_G262_,
    new_G267_, new_G268_, new_G269_, new_G3475_, new_G3482_, new_G2547_,
    new_G2554_, new_G386_, new_G389_, new_G392_, new_G395_, new_G1326_,
    new_G1329_, new_G1332_, new_G1436_, new_G1440_, new_G1445_, new_G1450_,
    new_G1454_, new_G2859_, new_G4385_, new_G3148_, new_G3239_, new_G3240_,
    new_G3265_, new_G3267_, new_G3270_, new_G3274_, new_G3277_, new_G3613_,
    new_G4515_, new_G4959_, new_G5000_, new_G5029_, new_G5117_, new_G5599_,
    new_G5687_, new_G6066_, new_G6124_, new_G6182_, new_G6934_, new_G6992_,
    new_G375_, new_G378_, new_G381_, new_G384_, new_G1328_, new_G1331_,
    new_G1334_, new_G1447_, new_G1766_, new_G2571_, new_G2579_, new_G2812_,
    new_G2816_, new_G2851_, new_G2861_, new_G6355_, new_G2863_, new_G6365_,
    new_G2866_, new_G3147_, new_G3242_, new_G3271_, new_G3279_, new_G3615_,
    new_G6843_, new_G3617_, new_G6851_, new_G3620_, new_G4056_, new_G4517_,
    new_G7451_, new_G4519_, new_G7461_, new_G4522_, new_G5031_, new_G5119_,
    new_G5481_, new_G5484_, new_G5539_, new_G5542_, new_G5601_, new_G5689_,
    new_G6067_, new_G6125_, new_G6183_, new_G6277_, new_G6280_, new_G6935_,
    new_G6993_, new_G7057_, new_G7060_, new_G7145_, new_G7148_, new_G4968_,
    new_G5009_, new_G2850_, new_G2862_, new_G2865_, new_G3149_, new_G3243_,
    new_G3616_, new_G3619_, new_G4518_, new_G4521_, new_G4965_, new_G5006_,
    new_G5483_, new_G5541_, new_G6279_, new_G7059_, new_G7147_, new_G374_,
    new_G377_, new_G380_, new_G383_, new_G955_, new_G4967_, new_G5008_,
    new_G975_, new_G1136_, new_G1140_, new_G1143_, new_G1145_, new_G1160_,
    new_G1771_, new_G1964_, new_G1968_, new_G1971_, new_G1973_, new_G2007_,
    new_G2578_, new_G2864_, new_G2867_, new_G3150_, new_G3245_, new_G3618_,
    new_G3621_, new_G4067_, new_G4520_, new_G4523_, new_G4713_, new_G4753_,
    new_G5037_, new_G5040_, new_G5125_, new_G5128_, new_G5485_, new_G5543_,
    new_G5607_, new_G5610_, new_G5695_, new_G5698_, new_G6073_, new_G6076_,
    new_G6131_, new_G6134_, new_G6189_, new_G6192_, new_G6281_, new_G6941_,
    new_G6944_, new_G6999_, new_G7002_, new_G7061_, new_G7149_, new_G958_,
    new_G967_, new_G971_, new_G1161_, new_G2008_, new_G2580_, new_G2868_,
    new_G3152_, new_G4443_, new_G4524_, new_G4721_, new_G4729_, new_G4737_,
    new_G4745_, new_G4761_, new_G4769_, new_G4777_, new_G4785_, new_G5039_,
    new_G5127_, new_G5609_, new_G5697_, new_G6075_, new_G6133_, new_G6191_,
    new_G6943_, new_G7001_, new_G3248_, new_G248_, new_G4719_, new_G294_,
    new_G4759_, new_G323_, new_G980_, new_G4072_, new_G5041_, new_G5129_,
    new_G5491_, new_G5494_, new_G5549_, new_G5552_, new_G5611_, new_G5699_,
    new_G6077_, new_G6135_, new_G6193_, new_G6287_, new_G6290_, new_G6945_,
    new_G7003_, new_G7067_, new_G7070_, new_G7155_, new_G7158_, new_G247_,
    new_G3155_, new_G251_, new_G272_, new_G961_, new_G275_, new_G293_,
    new_G297_, new_G300_, new_G303_, new_G306_, new_G4727_, new_G309_,
    new_G4735_, new_G312_, new_G4743_, new_G315_, new_G4751_, new_G318_,
    new_G322_, new_G4767_, new_G326_, new_G4775_, new_G329_, new_G4783_,
    new_G332_, new_G4791_, new_G335_, new_G2881_, new_G993_, new_G994_,
    new_G1166_, new_G1171_, new_G1174_, new_G2014_, new_G3459_, new_G3462_,
    new_G3464_, new_G3465_, new_G3490_, new_G4793_, new_G5493_, new_G5551_,
    new_G6289_, new_G7069_, new_G7157_, new_G250_, new_G274_, new_G308_,
    new_G311_, new_G314_, new_G317_, new_G325_, new_G328_, new_G331_,
    new_G334_, new_G417_, new_G991_, new_G992_, new_G3491_, new_G4801_,
    new_G4809_, new_G4817_, new_G4825_, new_G5047_, new_G5050_, new_G5135_,
    new_G5138_, new_G5495_, new_G5553_, new_G5617_, new_G5620_, new_G5705_,
    new_G5708_, new_G6083_, new_G6086_, new_G6141_, new_G6144_, new_G6199_,
    new_G6202_, new_G6291_, new_G6951_, new_G6954_, new_G7009_, new_G7012_,
    new_G7071_, new_G7159_, new_G271_, new_G296_, new_G299_, new_G302_,
    new_G305_, new_G4799_, new_G343_, new_G1170_, new_G1173_, new_G5049_,
    new_G5137_, new_G5167_, new_G5619_, new_G5707_, new_G6085_, new_G6143_,
    new_G6201_, new_G6953_, new_G7011_, new_G342_, new_G346_, new_G349_,
    new_G352_, new_G355_, new_G4807_, new_G358_, new_G4815_, new_G361_,
    new_G4823_, new_G364_, new_G4831_, new_G367_, new_G1172_, new_G1175_,
    new_G3497_, new_G5051_, new_G5139_, new_G5501_, new_G5504_, new_G5559_,
    new_G5562_, new_G5621_, new_G5709_, new_G6087_, new_G6145_, new_G6203_,
    new_G6297_, new_G6300_, new_G6955_, new_G7013_, new_G7077_, new_G7080_,
    new_G7165_, new_G7168_, new_G357_, new_G360_, new_G363_, new_G366_,
    new_G5173_, new_G5503_, new_G5561_, new_G6299_, new_G7079_, new_G7167_,
    new_G345_, new_G348_, new_G351_, new_G354_, new_G5057_, new_G5060_,
    new_G5145_, new_G5148_, new_G5505_, new_G5563_, new_G5627_, new_G5630_,
    new_G5715_, new_G5718_, new_G6093_, new_G6096_, new_G6151_, new_G6154_,
    new_G6209_, new_G6212_, new_G6301_, new_G6961_, new_G6964_, new_G7019_,
    new_G7022_, new_G7081_, new_G7169_, new_G5059_, new_G5147_, new_G5629_,
    new_G5717_, new_G6095_, new_G6153_, new_G6211_, new_G6963_, new_G7021_,
    new_G5061_, new_G5149_, new_G5511_, new_G5514_, new_G5569_, new_G5572_,
    new_G5631_, new_G5719_, new_G6097_, new_G6155_, new_G6213_, new_G6307_,
    new_G6310_, new_G6965_, new_G7023_, new_G7087_, new_G7090_, new_G7175_,
    new_G7178_, new_G5513_, new_G5571_, new_G6309_, new_G7089_, new_G7177_,
    new_G5067_, new_G5070_, new_G5155_, new_G5158_, new_G5515_, new_G5573_,
    new_G5637_, new_G5640_, new_G5725_, new_G5728_, new_G6103_, new_G6106_,
    new_G6161_, new_G6164_, new_G6219_, new_G6222_, new_G6311_, new_G6971_,
    new_G6974_, new_G7029_, new_G7032_, new_G7091_, new_G7179_, new_G5069_,
    new_G5157_, new_G5639_, new_G5727_, new_G6105_, new_G6163_, new_G6221_,
    new_G6973_, new_G7031_, new_G5521_, new_G1756_, new_G5579_, new_G1761_,
    new_G5071_, new_G5159_, new_G5641_, new_G5729_, new_G6107_, new_G6165_,
    new_G6223_, new_G6317_, new_G6320_, new_G6975_, new_G7033_, new_G7097_,
    new_G7100_, new_G7185_, new_G7188_, new_G1755_, new_G1760_, new_G6319_,
    new_G7099_, new_G7187_, new_G1757_, new_G1762_, new_G6113_, new_G2818_,
    new_G6171_, new_G2823_, new_G6981_, new_G4058_, new_G7039_, new_G4063_,
    new_G5077_, new_G5080_, new_G5165_, new_G5090_, new_G5647_, new_G5650_,
    new_G5735_, new_G5660_, new_G6229_, new_G6232_, new_G6321_, new_G7101_,
    new_G7189_, new_G2817_, new_G2822_, new_G4057_, new_G4062_, new_G5079_,
    new_G5089_, new_G5649_, new_G5659_, new_G6231_, new_G1782_, new_G1783_,
    new_G1784_, new_G1785_, new_G2819_, new_G2824_, new_G4059_, new_G4064_,
    new_G5081_, new_G5091_, new_G5651_, new_G5661_, new_G6233_, new_G6327_,
    new_G6252_, new_G7107_, new_G7110_, new_G7195_, new_G7120_, new_G5737_,
    new_G6251_, new_G7109_, new_G7119_, new_G5087_, new_G985_, new_G5097_,
    new_G988_, new_G5657_, new_G1776_, new_G5667_, new_G1779_, new_G2844_,
    new_G2845_, new_G2846_, new_G2847_, new_G4083_, new_G4084_, new_G4085_,
    new_G4086_, new_G6239_, new_G6242_, new_G6253_, new_G7111_, new_G7121_,
    new_G984_, new_G987_, new_G1775_, new_G1778_, new_G5743_, new_G6241_,
    new_G6329_, new_G7197_, new_G986_, new_G989_, new_G1777_, new_G1780_,
    new_G6259_, new_G2841_, new_G7117_, new_G4077_, new_G7127_, new_G4080_,
    new_G6243_, new_G990_, new_G996_, new_G1781_, new_G1787_, new_G2840_,
    new_G6335_, new_G4076_, new_G4079_, new_G7203_, new_G995_, new_G1786_,
    new_G6249_, new_G2838_, new_G2842_, new_G4078_, new_G4081_, new_G2837_,
    new_G2843_, new_G4082_, new_G4088_, new_G5170_, new_G5740_, new_G2839_,
    new_G2848_, new_G4087_, new_G1791_, new_G1003_, new_G5174_, new_G5744_,
    new_G2849_, new_G7200_, new_G1792_, new_G1004_, new_G6332_, new_G320_,
    new_G337_, new_G4092_, new_G7204_, new_G4093_, new_G2855_, new_G6336_,
    new_G369_, new_G2856_, new_G398_;
  assign G2 = G1;
  assign G3 = G1;
  assign new_G400_ = ~G57;
  assign new_G1184_ = G134 & G133;
  assign G450 = G1459;
  assign G448 = G1469;
  assign G444 = G1480;
  assign G442 = G1486;
  assign G440 = G1492;
  assign G438 = G1496;
  assign new_G1501_ = G199 & G188 & G162 & G172;
  assign G496 = G2208;
  assign G494 = G2218;
  assign G492 = G2224;
  assign G490 = G2230;
  assign G488 = G2236;
  assign G486 = G2239;
  assign G484 = G2247;
  assign G482 = G2253;
  assign G480 = G2256;
  assign new_G2857_ = G240 & G228 & G150 & G184;
  assign G560 = G3698;
  assign G542 = G3701;
  assign G558 = G3705;
  assign G556 = G3711;
  assign G554 = G3717;
  assign G552 = G3723;
  assign G550 = G3729;
  assign G548 = G3737;
  assign G546 = G3743;
  assign G544 = G3749;
  assign G540 = G4393;
  assign G538 = G4400;
  assign G536 = G4405;
  assign G534 = G4410;
  assign G532 = G4415;
  assign G530 = G4420;
  assign G528 = G4427;
  assign G526 = G4432;
  assign G524 = G4437;
  assign new_G4442_ = G186 & G185 & G183 & G182;
  assign new_G4514_ = G230 & G218 & G210 & G152;
  assign G279 = ~G15;
  assign new_G401_ = ~G5;
  assign new_G573_ = G1;
  assign new_G574_ = ~G5;
  assign new_G575_ = ~G5;
  assign new_G1178_ = ~G2236;
  assign new_G1186_ = ~G2253;
  assign new_G1192_ = ~G2256;
  assign new_G1198_ = G38;
  assign new_G1205_ = G15;
  assign new_G1206_ = ~G12 | ~G9;
  assign new_G1207_ = ~G12 | ~G9;
  assign new_G1210_ = G38;
  assign new_G1458_ = ~G1455;
  assign new_G1461_ = ~G1459;
  assign G436 = G1462;
  assign new_G1464_ = ~G1462;
  assign new_G1471_ = ~G1469;
  assign new_G1475_ = G106;
  assign new_G1482_ = ~G1480;
  assign new_G1488_ = ~G1486;
  assign new_G1495_ = ~G1492;
  assign new_G1499_ = ~G1496;
  assign new_G1500_ = ~G106;
  assign new_G1503_ = G18;
  assign new_G1512_ = G18;
  assign new_G1518_ = G4528 & G1492;
  assign new_G1524_ = G18;
  assign new_G1535_ = ~G18;
  assign new_G1541_ = ~G4528 | ~G1496;
  assign new_G2207_ = ~G2204;
  assign new_G2210_ = ~G2208;
  assign G478 = G2211;
  assign new_G2213_ = ~G2211;
  assign new_G2220_ = ~G2218;
  assign new_G2226_ = ~G2224;
  assign new_G2232_ = ~G2230;
  assign new_G2238_ = ~G2236;
  assign new_G2241_ = ~G2239;
  assign new_G2249_ = ~G2247;
  assign new_G2255_ = ~G2253;
  assign new_G2258_ = ~G2256;
  assign new_G2828_ = G4526;
  assign new_G3700_ = ~G3698;
  assign new_G3703_ = ~G3701;
  assign new_G3707_ = ~G3705;
  assign new_G3713_ = ~G3711;
  assign new_G3719_ = ~G3717;
  assign new_G3725_ = ~G3723;
  assign new_G3731_ = ~G3729;
  assign new_G3739_ = ~G3737;
  assign new_G3745_ = ~G3743;
  assign new_G3751_ = ~G3749;
  assign new_G4121_ = ~G4393;
  assign G522 = G4394;
  assign new_G4396_ = ~G4394;
  assign new_G4402_ = ~G4400;
  assign new_G4407_ = ~G4405;
  assign new_G4412_ = ~G4410;
  assign new_G4417_ = ~G4415;
  assign new_G4422_ = ~G4420;
  assign new_G4429_ = ~G4427;
  assign new_G4434_ = ~G4432;
  assign new_G4439_ = ~G4437;
  assign new_G4833_ = G4526;
  assign G402 = ~new_G400_ | ~new_G401_;
  assign G404 = ~new_G2857_;
  assign G406 = ~new_G4514_;
  assign G408 = ~new_G4442_;
  assign G410 = ~new_G1501_;
  assign new_G2876_ = new_G2857_ & new_G4514_;
  assign new_G2878_ = new_G4442_ & new_G1501_;
  assign G432 = new_G573_;
  assign G446 = new_G1475_;
  assign new_G1519_ = ~new_G1518_;
  assign new_G2871_ = G4528 & new_G1458_;
  assign new_G2883_ = ~G4528 | ~new_G2207_;
  assign new_G280_ = new_G1184_ & new_G575_;
  assign G284 = ~G1197 | ~new_G574_;
  assign G286 = ~new_G1205_;
  assign G289 = ~G1197 | ~new_G574_;
  assign G292 = ~new_G1184_ | ~new_G575_;
  assign G341 = ~new_G1205_;
  assign new_G4839_ = ~new_G4833_;
  assign new_G572_ = new_G573_;
  assign new_G581_ = new_G1206_;
  assign new_G587_ = new_G1512_;
  assign new_G601_ = new_G1206_;
  assign new_G606_ = new_G1512_;
  assign new_G650_ = new_G1206_;
  assign new_G657_ = new_G1512_;
  assign new_G671_ = new_G1207_;
  assign new_G678_ = new_G1503_;
  assign new_G777_ = new_G1541_ & new_G1198_;
  assign new_G1115_ = new_G1541_ & new_G1198_;
  assign new_G1336_ = new_G1512_;
  assign new_G1350_ = new_G1503_;
  assign new_G1477_ = ~new_G1475_;
  assign new_G1507_ = ~new_G1503_;
  assign new_G1514_ = ~new_G1512_;
  assign new_G1530_ = ~new_G1524_;
  assign new_G2259_ = new_G1535_;
  assign new_G2833_ = ~new_G2828_;
  assign new_G2872_ = ~new_G2871_;
  assign new_G2886_ = new_G1207_;
  assign new_G2892_ = new_G1503_;
  assign new_G2905_ = new_G1207_;
  assign new_G2909_ = new_G1503_;
  assign new_G3622_ = new_G1524_;
  assign new_G3635_ = new_G1524_;
  assign new_G3755_ = new_G1535_;
  assign new_G4640_ = new_G1524_;
  assign new_G4653_ = new_G1524_;
  assign new_G4873_ = new_G1541_;
  assign new_G4876_ = new_G1198_;
  assign new_G4881_ = new_G1488_;
  assign new_G4889_ = new_G1482_;
  assign new_G4905_ = new_G1471_;
  assign new_G4916_ = new_G1198_;
  assign new_G4921_ = new_G1464_;
  assign new_G5175_ = new_G1541_;
  assign new_G5178_ = new_G1198_;
  assign new_G5186_ = new_G1198_;
  assign new_G5191_ = new_G1488_;
  assign new_G5199_ = new_G1482_;
  assign new_G5215_ = new_G1471_;
  assign new_G5223_ = new_G1464_;
  assign new_G5393_ = new_G1192_;
  assign new_G5401_ = new_G1186_;
  assign new_G5409_ = new_G2249_;
  assign new_G5417_ = new_G1178_;
  assign new_G5425_ = new_G2232_;
  assign new_G5433_ = new_G2226_;
  assign new_G5441_ = new_G2220_;
  assign new_G5449_ = new_G2241_;
  assign new_G5457_ = new_G2213_;
  assign new_G5745_ = new_G1192_;
  assign new_G5753_ = new_G1186_;
  assign new_G5761_ = new_G2249_;
  assign new_G5769_ = new_G2241_;
  assign new_G5777_ = new_G1178_;
  assign new_G5785_ = new_G2232_;
  assign new_G5793_ = new_G2226_;
  assign new_G5801_ = new_G2220_;
  assign new_G5809_ = new_G2213_;
  assign new_G5865_ = new_G3751_;
  assign new_G5873_ = new_G3745_;
  assign new_G5881_ = new_G3739_;
  assign new_G5889_ = new_G3731_;
  assign new_G5897_ = new_G3725_;
  assign new_G5905_ = new_G3719_;
  assign new_G5913_ = new_G3713_;
  assign new_G5921_ = new_G3707_;
  assign new_G5985_ = new_G3751_;
  assign new_G5993_ = new_G3745_;
  assign new_G6001_ = new_G3739_;
  assign new_G6009_ = new_G3725_;
  assign new_G6017_ = new_G3719_;
  assign new_G6025_ = new_G3713_;
  assign new_G6033_ = new_G3707_;
  assign new_G6041_ = new_G3731_;
  assign new_G6514_ = new_G1210_;
  assign new_G6554_ = new_G1210_;
  assign new_G6567_ = new_G4439_;
  assign new_G6575_ = new_G4434_;
  assign new_G6583_ = new_G4429_;
  assign new_G6591_ = new_G4422_;
  assign new_G6599_ = new_G4417_;
  assign new_G6607_ = new_G4412_;
  assign new_G6615_ = new_G4407_;
  assign new_G6623_ = new_G4402_;
  assign new_G6631_ = new_G4396_;
  assign new_G6853_ = new_G4439_;
  assign new_G6861_ = new_G4434_;
  assign new_G6869_ = new_G4429_;
  assign new_G6877_ = new_G4417_;
  assign new_G6885_ = new_G4412_;
  assign new_G6893_ = new_G4407_;
  assign new_G6901_ = new_G4402_;
  assign new_G6909_ = new_G4422_;
  assign new_G6917_ = new_G4396_;
  assign G281 = ~new_G280_;
  assign G453 = new_G572_;
  assign new_G784_ = new_G1519_ & new_G1198_;
  assign new_G1014_ = new_G1198_ & new_G1519_;
  assign new_G3221_ = new_G2883_ & new_G1210_;
  assign new_G4913_ = new_G1519_;
  assign new_G4929_ = ~new_G1519_ & ~new_G1198_;
  assign new_G5183_ = new_G1519_;
  assign new_G5231_ = ~new_G1198_ & ~new_G1519_;
  assign new_G6511_ = new_G2883_;
  assign G278 = G163 & new_G572_;
  assign new_G615_ = G170 & new_G587_;
  assign new_G594_ = ~new_G587_;
  assign new_G611_ = ~new_G606_;
  assign new_G617_ = G169 & new_G587_;
  assign new_G619_ = G168 & new_G587_;
  assign new_G621_ = G167 & new_G587_;
  assign new_G623_ = G166 & new_G606_;
  assign new_G625_ = G165 & new_G606_;
  assign new_G627_ = G164 & new_G606_;
  assign new_G664_ = ~new_G657_;
  assign new_G685_ = ~new_G678_;
  assign new_G691_ = G177 & new_G657_;
  assign new_G693_ = G176 & new_G657_;
  assign new_G695_ = G175 & new_G657_;
  assign new_G697_ = G174 & new_G657_;
  assign new_G699_ = G173 & new_G657_;
  assign new_G701_ = G157 & new_G678_;
  assign new_G703_ = G156 & new_G678_;
  assign new_G705_ = G155 & new_G678_;
  assign new_G707_ = G154 & new_G678_;
  assign new_G709_ = G153 & new_G678_;
  assign new_G4879_ = ~new_G4873_;
  assign new_G4880_ = ~new_G4876_;
  assign new_G4887_ = ~new_G4881_;
  assign new_G4895_ = ~new_G4889_;
  assign new_G4911_ = ~new_G4905_;
  assign new_G4920_ = ~new_G4916_;
  assign new_G4927_ = ~new_G4921_;
  assign new_G5181_ = ~new_G5175_;
  assign new_G5182_ = ~new_G5178_;
  assign new_G5190_ = ~new_G5186_;
  assign new_G5197_ = ~new_G5191_;
  assign new_G5205_ = ~new_G5199_;
  assign new_G5221_ = ~new_G5215_;
  assign new_G5229_ = ~new_G5223_;
  assign new_G1343_ = ~new_G1336_;
  assign new_G1357_ = ~new_G1350_;
  assign new_G1364_ = G181 & new_G1336_;
  assign new_G1366_ = G171 & new_G1336_;
  assign new_G1368_ = G180 & new_G1336_;
  assign new_G1370_ = G179 & new_G1336_;
  assign new_G1372_ = G178 & new_G1336_;
  assign new_G1374_ = G161 & new_G1350_;
  assign new_G1376_ = G151 & new_G1350_;
  assign new_G1378_ = G160 & new_G1350_;
  assign new_G1380_ = G159 & new_G1350_;
  assign new_G1382_ = G158 & new_G1350_;
  assign new_G5399_ = ~new_G5393_;
  assign new_G5407_ = ~new_G5401_;
  assign new_G5415_ = ~new_G5409_;
  assign new_G5423_ = ~new_G5417_;
  assign new_G5431_ = ~new_G5425_;
  assign new_G5439_ = ~new_G5433_;
  assign new_G5447_ = ~new_G5441_;
  assign new_G5455_ = ~new_G5449_;
  assign new_G5463_ = ~new_G5457_;
  assign new_G5751_ = ~new_G5745_;
  assign new_G5759_ = ~new_G5753_;
  assign new_G5767_ = ~new_G5761_;
  assign new_G5775_ = ~new_G5769_;
  assign new_G5783_ = ~new_G5777_;
  assign new_G5791_ = ~new_G5785_;
  assign new_G5799_ = ~new_G5793_;
  assign new_G5807_ = ~new_G5801_;
  assign new_G5815_ = ~new_G5809_;
  assign new_G2019_ = new_G1514_;
  assign new_G2032_ = new_G1507_;
  assign new_G2117_ = new_G1514_;
  assign new_G2130_ = new_G1507_;
  assign new_G2266_ = ~new_G2259_;
  assign new_G2272_ = new_G1507_;
  assign new_G2286_ = G44 & new_G2259_;
  assign new_G2288_ = G41 & new_G2259_;
  assign new_G2290_ = G29 & new_G2259_;
  assign new_G2292_ = G26 & new_G2259_;
  assign new_G2294_ = G23 & new_G2259_;
  assign new_G5871_ = ~new_G5865_;
  assign new_G5879_ = ~new_G5873_;
  assign new_G5887_ = ~new_G5881_;
  assign new_G5895_ = ~new_G5889_;
  assign new_G5903_ = ~new_G5897_;
  assign new_G5911_ = ~new_G5905_;
  assign new_G5919_ = ~new_G5913_;
  assign new_G5927_ = ~new_G5921_;
  assign new_G5991_ = ~new_G5985_;
  assign new_G5999_ = ~new_G5993_;
  assign new_G6007_ = ~new_G6001_;
  assign new_G6015_ = ~new_G6009_;
  assign new_G6023_ = ~new_G6017_;
  assign new_G6031_ = ~new_G6025_;
  assign new_G6039_ = ~new_G6033_;
  assign new_G6047_ = ~new_G6041_;
  assign new_G2899_ = ~new_G2892_;
  assign new_G2914_ = ~new_G2909_;
  assign new_G2919_ = G209 & new_G2892_;
  assign new_G2921_ = G216 & new_G2892_;
  assign new_G2923_ = G215 & new_G2892_;
  assign new_G2925_ = G214 & new_G2892_;
  assign new_G2927_ = G213 & new_G2909_;
  assign new_G2929_ = G212 & new_G2909_;
  assign new_G2931_ = G211 & new_G2909_;
  assign new_G6518_ = ~new_G6514_;
  assign new_G3173_ = new_G2872_ & new_G1210_;
  assign new_G6558_ = ~new_G6554_;
  assign new_G6573_ = ~new_G6567_;
  assign new_G6581_ = ~new_G6575_;
  assign new_G6589_ = ~new_G6583_;
  assign new_G6597_ = ~new_G6591_;
  assign new_G6605_ = ~new_G6599_;
  assign new_G6613_ = ~new_G6607_;
  assign new_G6621_ = ~new_G6615_;
  assign new_G6629_ = ~new_G6623_;
  assign new_G6637_ = ~new_G6631_;
  assign new_G3629_ = ~new_G3622_;
  assign new_G3642_ = ~new_G3635_;
  assign new_G3649_ = new_G1461_ & new_G3622_;
  assign new_G3651_ = new_G1464_ & new_G3622_;
  assign new_G3653_ = new_G1471_ & new_G3622_;
  assign new_G3655_ = new_G1500_ & new_G3622_;
  assign new_G3657_ = new_G1482_ & new_G3622_;
  assign new_G3659_ = new_G1488_ & new_G3635_;
  assign new_G3661_ = new_G1495_ & new_G3635_;
  assign new_G3663_ = new_G1499_ & new_G3635_;
  assign new_G3762_ = ~new_G3755_;
  assign new_G3768_ = new_G1507_;
  assign new_G3782_ = G47 & new_G3755_;
  assign new_G3784_ = G35 & new_G3755_;
  assign new_G3786_ = G32 & new_G3755_;
  assign new_G3788_ = G50 & new_G3755_;
  assign new_G3790_ = G66 & new_G3755_;
  assign new_G6859_ = ~new_G6853_;
  assign new_G6867_ = ~new_G6861_;
  assign new_G6875_ = ~new_G6869_;
  assign new_G6883_ = ~new_G6877_;
  assign new_G6891_ = ~new_G6885_;
  assign new_G6899_ = ~new_G6893_;
  assign new_G6907_ = ~new_G6901_;
  assign new_G6915_ = ~new_G6909_;
  assign new_G6923_ = ~new_G6917_;
  assign new_G4094_ = new_G1530_;
  assign new_G4107_ = new_G1530_;
  assign new_G4444_ = new_G1530_;
  assign new_G4457_ = new_G1530_;
  assign new_G4647_ = ~new_G4640_;
  assign new_G4660_ = ~new_G4653_;
  assign new_G4667_ = new_G2210_ & new_G4640_;
  assign new_G4669_ = new_G2213_ & new_G4640_;
  assign new_G4671_ = new_G2220_ & new_G4640_;
  assign new_G4673_ = new_G2226_ & new_G4640_;
  assign new_G4675_ = new_G2232_ & new_G4640_;
  assign new_G4677_ = new_G2238_ & new_G4653_;
  assign new_G4679_ = new_G2241_ & new_G4653_;
  assign new_G4681_ = new_G2249_ & new_G4653_;
  assign new_G4683_ = new_G2255_ & new_G4653_;
  assign new_G4685_ = new_G2258_ & new_G4653_;
  assign new_G4897_ = new_G1477_;
  assign new_G5207_ = new_G1477_;
  assign new_G6551_ = new_G2872_;
  assign new_G763_ = ~new_G4876_ | ~new_G4879_;
  assign new_G764_ = ~new_G4873_ | ~new_G4880_;
  assign new_G4919_ = ~new_G4913_;
  assign new_G886_ = ~new_G4913_ | ~new_G4920_;
  assign new_G1005_ = ~new_G5178_ | ~new_G5181_;
  assign new_G1006_ = ~new_G5175_ | ~new_G5182_;
  assign new_G5189_ = ~new_G5183_;
  assign new_G1018_ = ~new_G5183_ | ~new_G5190_;
  assign new_G5237_ = ~new_G5231_;
  assign new_G6517_ = ~new_G6511_;
  assign new_G3169_ = ~new_G6511_ | ~new_G6518_;
  assign new_G4935_ = ~new_G4929_;
  assign new_G4970_ = new_G784_;
  assign new_G5239_ = new_G1014_;
  assign new_G577_ = new_G594_ | new_G615_;
  assign new_G616_ = new_G594_ | new_G587_;
  assign new_G618_ = new_G594_ | new_G617_;
  assign new_G620_ = new_G594_ | new_G619_;
  assign new_G622_ = new_G594_ | new_G621_;
  assign new_G624_ = new_G611_ | new_G623_;
  assign new_G626_ = new_G611_ | new_G625_;
  assign new_G628_ = new_G611_ | new_G627_;
  assign new_G692_ = new_G664_ | new_G691_;
  assign new_G694_ = new_G664_ | new_G693_;
  assign new_G696_ = new_G664_ | new_G695_;
  assign new_G698_ = new_G664_ | new_G697_;
  assign new_G700_ = new_G664_ | new_G699_;
  assign new_G702_ = new_G685_ | new_G701_;
  assign new_G704_ = new_G685_ | new_G703_;
  assign new_G706_ = new_G685_ | new_G705_;
  assign new_G708_ = new_G685_ | new_G707_;
  assign new_G710_ = new_G685_ | new_G709_;
  assign new_G765_ = ~new_G763_ | ~new_G764_;
  assign new_G4903_ = ~new_G4897_;
  assign new_G885_ = ~new_G4916_ | ~new_G4919_;
  assign new_G1007_ = ~new_G1005_ | ~new_G1006_;
  assign new_G1017_ = ~new_G5186_ | ~new_G5189_;
  assign new_G5213_ = ~new_G5207_;
  assign new_G1363_ = G141 & new_G1343_;
  assign new_G1365_ = G147 & new_G1343_;
  assign new_G1367_ = G138 & new_G1343_;
  assign new_G1369_ = G144 & new_G1343_;
  assign new_G1371_ = G135 & new_G1343_;
  assign new_G1373_ = G141 & new_G1357_;
  assign new_G1375_ = G147 & new_G1357_;
  assign new_G1377_ = G138 & new_G1357_;
  assign new_G1379_ = G144 & new_G1357_;
  assign new_G1381_ = G135 & new_G1357_;
  assign new_G2026_ = ~new_G2019_;
  assign new_G2039_ = ~new_G2032_;
  assign new_G2046_ = G103 & new_G2019_;
  assign new_G2048_ = G130 & new_G2019_;
  assign new_G2050_ = G127 & new_G2019_;
  assign new_G2052_ = G124 & new_G2019_;
  assign new_G2054_ = G100 & new_G2019_;
  assign new_G2056_ = G103 & new_G2032_;
  assign new_G2058_ = G130 & new_G2032_;
  assign new_G2060_ = G127 & new_G2032_;
  assign new_G2062_ = G124 & new_G2032_;
  assign new_G2064_ = G100 & new_G2032_;
  assign new_G2124_ = ~new_G2117_;
  assign new_G2137_ = ~new_G2130_;
  assign new_G2144_ = G115 & new_G2117_;
  assign new_G2146_ = G118 & new_G2117_;
  assign new_G2148_ = G97 & new_G2117_;
  assign new_G2150_ = G94 & new_G2117_;
  assign new_G2152_ = G121 & new_G2117_;
  assign new_G2154_ = G115 & new_G2130_;
  assign new_G2156_ = G118 & new_G2130_;
  assign new_G2158_ = G97 & new_G2130_;
  assign new_G2160_ = G94 & new_G2130_;
  assign new_G2162_ = G121 & new_G2130_;
  assign new_G2279_ = ~new_G2272_;
  assign new_G2285_ = G208 & new_G2266_;
  assign new_G2287_ = G198 & new_G2266_;
  assign new_G2289_ = G207 & new_G2266_;
  assign new_G2291_ = G206 & new_G2266_;
  assign new_G2293_ = G205 & new_G2266_;
  assign new_G2296_ = G44 & new_G2272_;
  assign new_G2298_ = G41 & new_G2272_;
  assign new_G2300_ = G29 & new_G2272_;
  assign new_G2302_ = G26 & new_G2272_;
  assign new_G2304_ = G23 & new_G2272_;
  assign new_G2918_ = new_G2899_ | new_G2892_;
  assign new_G2920_ = new_G2899_ | new_G2919_;
  assign new_G2922_ = new_G2899_ | new_G2921_;
  assign new_G2924_ = new_G2899_ | new_G2923_;
  assign new_G2926_ = new_G2899_ | new_G2925_;
  assign new_G2928_ = new_G2914_ | new_G2927_;
  assign new_G2930_ = new_G2914_ | new_G2929_;
  assign new_G2932_ = new_G2914_ | new_G2931_;
  assign new_G3168_ = ~new_G6514_ | ~new_G6517_;
  assign new_G6557_ = ~new_G6551_;
  assign new_G3211_ = ~new_G6551_ | ~new_G6558_;
  assign new_G3648_ = G114 & new_G3629_;
  assign new_G3650_ = G113 & new_G3629_;
  assign new_G3652_ = G111 & new_G3629_;
  assign new_G3654_ = G87 & new_G3629_;
  assign new_G3656_ = G112 & new_G3629_;
  assign new_G3658_ = G88 & new_G3642_;
  assign new_G3660_ = G1455 & new_G3642_;
  assign new_G3662_ = G2204 & new_G3642_;
  assign new_G3665_ = new_G3703_ & new_G3642_;
  assign new_G3666_ = G70 & new_G3642_;
  assign new_G3775_ = ~new_G3768_;
  assign new_G3781_ = G193 & new_G3762_;
  assign new_G3783_ = G192 & new_G3762_;
  assign new_G3785_ = G191 & new_G3762_;
  assign new_G3787_ = G190 & new_G3762_;
  assign new_G3789_ = G189 & new_G3762_;
  assign new_G3792_ = G47 & new_G3768_;
  assign new_G3794_ = G35 & new_G3768_;
  assign new_G3796_ = G32 & new_G3768_;
  assign new_G3798_ = G50 & new_G3768_;
  assign new_G3800_ = G66 & new_G3768_;
  assign new_G4101_ = ~new_G4094_;
  assign new_G4114_ = ~new_G4107_;
  assign new_G4123_ = G58 & new_G4094_;
  assign new_G4126_ = G77 & new_G4094_;
  assign new_G4129_ = G78 & new_G4094_;
  assign new_G4132_ = G59 & new_G4094_;
  assign new_G4135_ = G81 & new_G4094_;
  assign new_G4138_ = G80 & new_G4107_;
  assign new_G4141_ = G79 & new_G4107_;
  assign new_G4144_ = G60 & new_G4107_;
  assign new_G4147_ = G61 & new_G4107_;
  assign new_G4150_ = G62 & new_G4107_;
  assign new_G4451_ = ~new_G4444_;
  assign new_G4464_ = ~new_G4457_;
  assign new_G4471_ = G69 & new_G4444_;
  assign new_G4473_ = G70 & new_G4444_;
  assign new_G4475_ = G74 & new_G4444_;
  assign new_G4477_ = G76 & new_G4444_;
  assign new_G4479_ = G75 & new_G4444_;
  assign new_G4481_ = G73 & new_G4457_;
  assign new_G4483_ = G53 & new_G4457_;
  assign new_G4485_ = G54 & new_G4457_;
  assign new_G4487_ = G55 & new_G4457_;
  assign new_G4489_ = G56 & new_G4457_;
  assign new_G4666_ = G82 & new_G4647_;
  assign new_G4668_ = G65 & new_G4647_;
  assign new_G4670_ = G83 & new_G4647_;
  assign new_G4672_ = G84 & new_G4647_;
  assign new_G4674_ = G85 & new_G4647_;
  assign new_G4676_ = G64 & new_G4660_;
  assign new_G4678_ = G63 & new_G4660_;
  assign new_G4680_ = G86 & new_G4660_;
  assign new_G4682_ = G109 & new_G4660_;
  assign new_G4684_ = G110 & new_G4660_;
  assign new_G579_ = new_G577_ & new_G581_;
  assign new_G629_ = new_G616_ & new_G581_;
  assign new_G633_ = new_G618_ & new_G581_;
  assign new_G637_ = new_G620_ & new_G581_;
  assign new_G641_ = new_G622_ & new_G581_;
  assign new_G645_ = new_G624_ & new_G601_;
  assign new_G711_ = new_G692_ & new_G650_;
  assign new_G715_ = new_G694_ & new_G650_;
  assign new_G719_ = new_G696_ & new_G650_;
  assign new_G723_ = new_G698_ & new_G650_;
  assign new_G727_ = new_G700_ & new_G650_;
  assign new_G731_ = new_G702_ & new_G671_;
  assign new_G737_ = new_G704_ & new_G671_;
  assign new_G745_ = new_G706_ & new_G671_;
  assign new_G751_ = new_G708_ & new_G671_;
  assign new_G757_ = new_G710_ & new_G671_;
  assign new_G887_ = ~new_G885_ | ~new_G886_;
  assign new_G1019_ = ~new_G1017_ | ~new_G1018_;
  assign new_G5245_ = ~new_G5239_;
  assign new_G1383_ = new_G1365_ | new_G1366_;
  assign new_G1387_ = new_G1367_ | new_G1368_;
  assign new_G1391_ = new_G1369_ | new_G1370_;
  assign new_G1395_ = new_G1371_ | new_G1372_;
  assign new_G1399_ = new_G1375_ | new_G1376_;
  assign new_G1406_ = new_G1377_ | new_G1378_;
  assign new_G1412_ = new_G1379_ | new_G1380_;
  assign new_G1418_ = new_G1381_ | new_G1382_;
  assign new_G2305_ = new_G2287_ | new_G2288_;
  assign new_G2308_ = new_G2289_ | new_G2290_;
  assign new_G2312_ = new_G2291_ | new_G2292_;
  assign new_G2316_ = new_G2293_ | new_G2294_;
  assign new_G2933_ = new_G2920_ & new_G2886_;
  assign new_G2938_ = new_G2922_ & new_G2886_;
  assign new_G2942_ = new_G2924_ & new_G2886_;
  assign new_G2946_ = new_G2926_ & new_G2886_;
  assign new_G2950_ = new_G2928_ & new_G2905_;
  assign new_G3170_ = ~new_G3168_ | ~new_G3169_;
  assign new_G3210_ = ~new_G6554_ | ~new_G6557_;
  assign new_G3667_ = new_G3650_ | new_G3651_;
  assign new_G3670_ = new_G3652_ | new_G3653_;
  assign new_G3673_ = new_G3654_ | new_G3655_;
  assign new_G3676_ = new_G3656_ | new_G3657_;
  assign new_G3679_ = new_G3658_ | new_G3659_;
  assign new_G3682_ = new_G3665_ | new_G3635_;
  assign new_G3686_ = new_G3666_ | new_G3635_;
  assign new_G3801_ = new_G3781_ | new_G3782_;
  assign new_G3804_ = new_G3783_ | new_G3784_;
  assign new_G3807_ = new_G3785_ | new_G3786_;
  assign new_G3810_ = new_G3787_ | new_G3788_;
  assign new_G3813_ = new_G3789_ | new_G3790_;
  assign new_G4525_ = new_G2918_ & new_G2886_;
  assign new_G4686_ = new_G4668_ | new_G4669_;
  assign new_G4689_ = new_G4670_ | new_G4671_;
  assign new_G4692_ = new_G4672_ | new_G4673_;
  assign new_G4695_ = new_G4674_ | new_G4675_;
  assign new_G4698_ = new_G4676_ | new_G4677_;
  assign new_G4701_ = new_G4678_ | new_G4679_;
  assign new_G4704_ = new_G4680_ | new_G4681_;
  assign new_G4707_ = new_G4682_ | new_G4683_;
  assign new_G4710_ = new_G4684_ | new_G4685_;
  assign new_G4976_ = ~new_G4970_;
  assign new_G5271_ = new_G2932_ & new_G2905_;
  assign new_G5274_ = new_G2930_ & new_G2905_;
  assign new_G5305_ = new_G628_ & new_G601_;
  assign new_G5308_ = new_G626_ & new_G601_;
  assign new_G5318_ = new_G1373_ | new_G1374_;
  assign new_G6690_ = new_G3648_ | new_G3649_;
  assign new_G6711_ = new_G3662_ | new_G3663_;
  assign new_G6714_ = new_G3660_ | new_G3661_;
  assign new_G7252_ = new_G2285_ | new_G2286_;
  assign new_G7296_ = new_G1363_ | new_G1364_;
  assign new_G7466_ = new_G4666_ | new_G4667_;
  assign new_G907_ = new_G765_ & new_G784_;
  assign new_G913_ = new_G765_ & new_G784_;
  assign new_G915_ = new_G765_ & new_G784_;
  assign new_G916_ = new_G765_ & new_G784_;
  assign new_G1116_ = new_G1007_ & new_G1014_;
  assign new_G2045_ = G204 & new_G2026_;
  assign new_G2047_ = G203 & new_G2026_;
  assign new_G2049_ = G202 & new_G2026_;
  assign new_G2051_ = G201 & new_G2026_;
  assign new_G2053_ = G200 & new_G2026_;
  assign new_G2055_ = G235 & new_G2039_;
  assign new_G2057_ = G234 & new_G2039_;
  assign new_G2059_ = G233 & new_G2039_;
  assign new_G2061_ = G232 & new_G2039_;
  assign new_G2063_ = G231 & new_G2039_;
  assign new_G2143_ = G197 & new_G2124_;
  assign new_G2145_ = G187 & new_G2124_;
  assign new_G2147_ = G196 & new_G2124_;
  assign new_G2149_ = G195 & new_G2124_;
  assign new_G2151_ = G194 & new_G2124_;
  assign new_G2153_ = G227 & new_G2137_;
  assign new_G2155_ = G217 & new_G2137_;
  assign new_G2157_ = G226 & new_G2137_;
  assign new_G2159_ = G225 & new_G2137_;
  assign new_G2161_ = G224 & new_G2137_;
  assign new_G2295_ = G239 & new_G2279_;
  assign new_G2297_ = G229 & new_G2279_;
  assign new_G2299_ = G238 & new_G2279_;
  assign new_G2301_ = G237 & new_G2279_;
  assign new_G2303_ = G236 & new_G2279_;
  assign new_G3212_ = ~new_G3210_ | ~new_G3211_;
  assign new_G3791_ = G223 & new_G3775_;
  assign new_G3793_ = G222 & new_G3775_;
  assign new_G3795_ = G221 & new_G3775_;
  assign new_G3797_ = G220 & new_G3775_;
  assign new_G3799_ = G219 & new_G3775_;
  assign new_G4122_ = new_G4121_ & new_G4101_;
  assign new_G4125_ = new_G4396_ & new_G4101_;
  assign new_G4128_ = new_G4402_ & new_G4101_;
  assign new_G4131_ = new_G4407_ & new_G4101_;
  assign new_G4134_ = new_G4412_ & new_G4101_;
  assign new_G4137_ = new_G4417_ & new_G4114_;
  assign new_G4140_ = new_G4422_ & new_G4114_;
  assign new_G4143_ = new_G4429_ & new_G4114_;
  assign new_G4146_ = new_G4434_ & new_G4114_;
  assign new_G4149_ = new_G4439_ & new_G4114_;
  assign new_G4470_ = new_G3700_ & new_G4451_;
  assign new_G4472_ = new_G3703_ & new_G4451_;
  assign new_G4474_ = new_G3707_ & new_G4451_;
  assign new_G4476_ = new_G3713_ & new_G4451_;
  assign new_G4478_ = new_G3719_ & new_G4451_;
  assign new_G4480_ = new_G3725_ & new_G4464_;
  assign new_G4482_ = new_G3731_ & new_G4464_;
  assign new_G4484_ = new_G3739_ & new_G4464_;
  assign new_G4486_ = new_G3745_ & new_G4464_;
  assign new_G4488_ = new_G3751_ & new_G4464_;
  assign new_G4962_ = new_G765_;
  assign new_G5003_ = new_G765_;
  assign new_G5234_ = new_G1007_;
  assign new_G5242_ = new_G1007_;
  assign new_G5250_ = ~new_G4525_;
  assign new_G5284_ = ~new_G579_;
  assign new_G802_ = new_G1488_ & new_G2950_;
  assign new_G821_ = new_G1482_ & new_G2946_;
  assign new_G845_ = new_G1477_ & new_G2942_;
  assign new_G868_ = new_G1471_ & new_G2938_;
  assign new_G877_ = new_G1464_ & new_G2933_;
  assign new_G902_ = new_G887_ & new_G765_;
  assign new_G908_ = new_G777_ | new_G907_;
  assign new_G914_ = new_G887_ & new_G765_;
  assign new_G917_ = new_G777_ | new_G916_;
  assign new_G953_ = new_G887_ & new_G765_;
  assign new_G1023_ = ~new_G1019_;
  assign new_G1035_ = new_G1488_ & new_G2950_;
  assign new_G1050_ = new_G1482_ & new_G2946_;
  assign new_G1068_ = new_G1477_ & new_G2942_;
  assign new_G1086_ = new_G1471_ & new_G2938_;
  assign new_G1102_ = new_G1464_ & new_G2933_;
  assign new_G1108_ = new_G1019_ & new_G1007_;
  assign new_G1117_ = new_G1115_ | new_G1116_;
  assign new_G5322_ = ~new_G5318_;
  assign new_G1553_ = new_G1192_ & new_G757_;
  assign new_G1567_ = new_G1186_ & new_G751_;
  assign new_G1584_ = new_G2249_ & new_G745_;
  assign new_G1590_ = new_G2241_ & new_G737_;
  assign new_G1606_ = new_G1178_ & new_G731_;
  assign new_G1624_ = new_G2232_ & new_G1418_;
  assign new_G1647_ = new_G2226_ & new_G1412_;
  assign new_G1669_ = new_G2220_ & new_G1406_;
  assign new_G1677_ = new_G2213_ & new_G1399_;
  assign new_G1802_ = new_G1192_ & new_G757_;
  assign new_G1816_ = new_G1186_ & new_G751_;
  assign new_G1834_ = new_G2249_ & new_G745_;
  assign new_G1841_ = new_G737_ & new_G2241_;
  assign new_G1866_ = new_G1178_ & new_G731_;
  assign new_G1880_ = new_G2232_ & new_G1418_;
  assign new_G1897_ = new_G2226_ & new_G1412_;
  assign new_G1914_ = new_G2220_ & new_G1406_;
  assign new_G1929_ = new_G2213_ & new_G1399_;
  assign new_G2065_ = new_G2045_ | new_G2046_;
  assign new_G2069_ = new_G2047_ | new_G2048_;
  assign new_G2073_ = new_G2049_ | new_G2050_;
  assign new_G2077_ = new_G2051_ | new_G2052_;
  assign new_G2081_ = new_G2053_ | new_G2054_;
  assign new_G2085_ = new_G2055_ | new_G2056_;
  assign new_G2091_ = new_G2057_ | new_G2058_;
  assign new_G2099_ = new_G2059_ | new_G2060_;
  assign new_G2105_ = new_G2061_ | new_G2062_;
  assign new_G2111_ = new_G2063_ | new_G2064_;
  assign new_G2163_ = new_G2145_ | new_G2146_;
  assign new_G2167_ = new_G2147_ | new_G2148_;
  assign new_G2171_ = new_G2149_ | new_G2150_;
  assign new_G2175_ = new_G2151_ | new_G2152_;
  assign new_G2179_ = new_G2155_ | new_G2156_;
  assign new_G2186_ = new_G2157_ | new_G2158_;
  assign new_G2192_ = new_G2159_ | new_G2160_;
  assign new_G2198_ = new_G2161_ | new_G2162_;
  assign new_G2320_ = new_G2297_ | new_G2298_;
  assign new_G2323_ = new_G2299_ | new_G2300_;
  assign new_G2329_ = new_G2301_ | new_G2302_;
  assign new_G2335_ = new_G2303_ | new_G2304_;
  assign new_G2962_ = new_G4710_ & new_G727_;
  assign new_G2970_ = new_G4707_ & new_G723_;
  assign new_G2977_ = new_G4704_ & new_G719_;
  assign new_G2979_ = new_G4701_ & new_G715_;
  assign new_G2989_ = new_G4698_ & new_G711_;
  assign new_G2998_ = new_G4695_ & new_G1395_;
  assign new_G3006_ = new_G4692_ & new_G1391_;
  assign new_G3013_ = new_G4689_ & new_G1387_;
  assign new_G3015_ = new_G4686_ & new_G1383_;
  assign new_G3183_ = new_G3679_ & new_G645_;
  assign new_G3192_ = new_G3676_ & new_G641_;
  assign new_G3200_ = new_G3673_ & new_G637_;
  assign new_G3207_ = new_G3670_ & new_G633_;
  assign new_G3209_ = new_G3667_ & new_G629_;
  assign new_G3216_ = new_G3212_ & new_G3170_;
  assign new_G3222_ = new_G3170_ & new_G3173_;
  assign new_G6694_ = ~new_G6690_;
  assign new_G3695_ = new_G1535_ & new_G2305_;
  assign new_G3816_ = new_G3791_ | new_G3792_;
  assign new_G3821_ = new_G3793_ | new_G3794_;
  assign new_G3828_ = new_G3795_ | new_G3796_;
  assign new_G3833_ = new_G3797_ | new_G3798_;
  assign new_G3838_ = new_G3799_ | new_G3800_;
  assign new_G4151_ = new_G4125_ | new_G4126_;
  assign new_G4154_ = new_G4128_ | new_G4129_;
  assign new_G4157_ = new_G4131_ | new_G4132_;
  assign new_G4160_ = new_G4134_ | new_G4135_;
  assign new_G4163_ = new_G4137_ | new_G4138_;
  assign new_G4166_ = new_G4140_ | new_G4141_;
  assign new_G4169_ = new_G4143_ | new_G4144_;
  assign new_G4172_ = new_G4146_ | new_G4147_;
  assign new_G4175_ = new_G4149_ | new_G4150_;
  assign new_G7256_ = ~new_G7252_;
  assign new_G7300_ = ~new_G7296_;
  assign new_G4490_ = new_G4474_ | new_G4475_;
  assign new_G4493_ = new_G4476_ | new_G4477_;
  assign new_G4496_ = new_G4478_ | new_G4479_;
  assign new_G4499_ = new_G4480_ | new_G4481_;
  assign new_G4502_ = new_G4482_ | new_G4483_;
  assign new_G4505_ = new_G4484_ | new_G4485_;
  assign new_G4508_ = new_G4486_ | new_G4487_;
  assign new_G4511_ = new_G4488_ | new_G4489_;
  assign new_G7470_ = ~new_G7466_;
  assign new_G4884_ = new_G2950_;
  assign new_G4892_ = new_G2946_;
  assign new_G4900_ = new_G2942_;
  assign new_G4908_ = new_G2938_;
  assign new_G4924_ = new_G2933_;
  assign new_G4952_ = new_G887_;
  assign new_G4983_ = ~new_G777_ & ~new_G915_;
  assign new_G4993_ = new_G887_;
  assign new_G5011_ = ~new_G1464_ & ~new_G2933_;
  assign new_G5194_ = new_G2950_;
  assign new_G5202_ = new_G2946_;
  assign new_G5210_ = new_G2942_;
  assign new_G5218_ = new_G2938_;
  assign new_G5226_ = new_G2933_;
  assign new_G5247_ = new_G2933_;
  assign new_G5255_ = new_G2942_;
  assign new_G5258_ = new_G2938_;
  assign new_G5263_ = new_G2950_;
  assign new_G5266_ = new_G2946_;
  assign new_G5277_ = ~new_G5271_;
  assign new_G5278_ = ~new_G5274_;
  assign new_G5281_ = new_G629_;
  assign new_G5289_ = new_G637_;
  assign new_G5292_ = new_G633_;
  assign new_G5297_ = new_G645_;
  assign new_G5300_ = new_G641_;
  assign new_G5311_ = ~new_G5305_;
  assign new_G5312_ = ~new_G5308_;
  assign new_G5315_ = new_G1399_;
  assign new_G5323_ = new_G1412_;
  assign new_G5326_ = new_G1406_;
  assign new_G5331_ = new_G731_;
  assign new_G5334_ = new_G1418_;
  assign new_G5339_ = new_G745_;
  assign new_G5342_ = new_G737_;
  assign new_G5349_ = new_G757_;
  assign new_G5352_ = new_G751_;
  assign new_G5396_ = new_G757_;
  assign new_G5404_ = new_G751_;
  assign new_G5412_ = new_G745_;
  assign new_G5420_ = new_G731_;
  assign new_G5428_ = new_G1418_;
  assign new_G5436_ = new_G1412_;
  assign new_G5444_ = new_G1406_;
  assign new_G5452_ = new_G737_;
  assign new_G5460_ = new_G1399_;
  assign new_G5465_ = ~new_G2241_ & ~new_G737_;
  assign new_G5581_ = ~new_G2213_ & ~new_G1399_;
  assign new_G5748_ = new_G757_;
  assign new_G5756_ = new_G751_;
  assign new_G5764_ = new_G745_;
  assign new_G5772_ = new_G737_;
  assign new_G5780_ = new_G731_;
  assign new_G5788_ = new_G1418_;
  assign new_G5796_ = new_G1412_;
  assign new_G5804_ = new_G1406_;
  assign new_G5812_ = new_G1399_;
  assign new_G5849_ = ~new_G737_ & ~new_G2241_;
  assign new_G5929_ = new_G3682_;
  assign new_G6049_ = new_G3682_;
  assign new_G6367_ = new_G4710_;
  assign new_G6370_ = new_G727_;
  assign new_G6375_ = new_G4707_;
  assign new_G6378_ = new_G723_;
  assign new_G6383_ = new_G4704_;
  assign new_G6386_ = new_G719_;
  assign new_G6391_ = new_G4698_;
  assign new_G6394_ = new_G711_;
  assign new_G6399_ = new_G4695_;
  assign new_G6402_ = new_G1395_;
  assign new_G6407_ = new_G4692_;
  assign new_G6410_ = new_G1391_;
  assign new_G6415_ = new_G4689_;
  assign new_G6418_ = new_G1387_;
  assign new_G6423_ = new_G4701_;
  assign new_G6426_ = new_G715_;
  assign new_G6431_ = new_G4686_;
  assign new_G6434_ = new_G1383_;
  assign new_G6442_ = new_G3813_;
  assign new_G6450_ = new_G3810_;
  assign new_G6458_ = new_G3807_;
  assign new_G6466_ = new_G3801_;
  assign new_G6498_ = new_G3804_;
  assign new_G6519_ = new_G3679_;
  assign new_G6522_ = new_G645_;
  assign new_G6527_ = new_G3676_;
  assign new_G6530_ = new_G641_;
  assign new_G6535_ = new_G3673_;
  assign new_G6538_ = new_G637_;
  assign new_G6543_ = new_G3670_;
  assign new_G6546_ = new_G633_;
  assign new_G6559_ = new_G3667_;
  assign new_G6562_ = new_G629_;
  assign new_G6687_ = new_G3667_;
  assign new_G6695_ = new_G3673_;
  assign new_G6698_ = new_G3670_;
  assign new_G6703_ = new_G3679_;
  assign new_G6706_ = new_G3676_;
  assign new_G6717_ = ~new_G6711_;
  assign new_G6718_ = ~new_G6714_;
  assign new_G6724_ = new_G2153_ | new_G2154_;
  assign new_G6768_ = new_G2295_ | new_G2296_;
  assign new_G7208_ = new_G2143_ | new_G2144_;
  assign new_G7221_ = new_G3801_;
  assign new_G7229_ = new_G3807_;
  assign new_G7232_ = new_G3804_;
  assign new_G7239_ = new_G3813_;
  assign new_G7242_ = new_G3810_;
  assign new_G7249_ = new_G2305_;
  assign new_G7257_ = new_G2312_;
  assign new_G7260_ = new_G2308_;
  assign new_G7268_ = new_G2316_;
  assign new_G7293_ = new_G1383_;
  assign new_G7301_ = new_G1391_;
  assign new_G7304_ = new_G1387_;
  assign new_G7309_ = new_G711_;
  assign new_G7312_ = new_G1395_;
  assign new_G7317_ = new_G719_;
  assign new_G7320_ = new_G715_;
  assign new_G7327_ = new_G727_;
  assign new_G7330_ = new_G723_;
  assign new_G7396_ = new_G2316_;
  assign new_G7404_ = new_G2312_;
  assign new_G7412_ = new_G2308_;
  assign new_G7425_ = new_G3686_;
  assign new_G7463_ = new_G4686_;
  assign new_G7471_ = new_G4692_;
  assign new_G7474_ = new_G4689_;
  assign new_G7479_ = new_G4698_;
  assign new_G7482_ = new_G4695_;
  assign new_G7487_ = new_G4704_;
  assign new_G7490_ = new_G4701_;
  assign new_G7497_ = new_G4710_;
  assign new_G7500_ = new_G4707_;
  assign new_G7507_ = new_G4472_ | new_G4473_;
  assign new_G7510_ = new_G4470_ | new_G4471_;
  assign new_G7554_ = new_G4122_ | new_G4123_;
  assign new_G1152_ = ~new_G5234_ | ~new_G5237_;
  assign new_G5238_ = ~new_G5234_;
  assign new_G1156_ = ~new_G5242_ | ~new_G5245_;
  assign new_G5246_ = ~new_G5242_;
  assign new_G5254_ = ~new_G5250_;
  assign new_G5288_ = ~new_G5284_;
  assign new_G3223_ = new_G3221_ | new_G3222_;
  assign new_G4942_ = new_G914_ | new_G777_ | new_G913_;
  assign new_G4966_ = ~new_G4962_;
  assign new_G5007_ = ~new_G5003_;
  assign new_G5279_ = ~new_G5274_ | ~new_G5277_;
  assign new_G5280_ = ~new_G5271_ | ~new_G5278_;
  assign new_G5313_ = ~new_G5308_ | ~new_G5311_;
  assign new_G5314_ = ~new_G5305_ | ~new_G5312_;
  assign new_G6719_ = ~new_G6714_ | ~new_G6717_;
  assign new_G6720_ = ~new_G6711_ | ~new_G6718_;
  assign new_G790_ = ~new_G4884_ | ~new_G4887_;
  assign new_G4888_ = ~new_G4884_;
  assign new_G803_ = ~new_G4892_ | ~new_G4895_;
  assign new_G4896_ = ~new_G4892_;
  assign new_G825_ = ~new_G4900_ | ~new_G4903_;
  assign new_G4904_ = ~new_G4900_;
  assign new_G851_ = ~new_G4908_ | ~new_G4911_;
  assign new_G4912_ = ~new_G4908_;
  assign new_G893_ = ~new_G4924_ | ~new_G4927_;
  assign new_G4928_ = ~new_G4924_;
  assign new_G906_ = ~new_G902_;
  assign new_G912_ = ~new_G908_;
  assign new_G1024_ = ~new_G5194_ | ~new_G5197_;
  assign new_G5198_ = ~new_G5194_;
  assign new_G1036_ = ~new_G5202_ | ~new_G5205_;
  assign new_G5206_ = ~new_G5202_;
  assign new_G1053_ = ~new_G5210_ | ~new_G5213_;
  assign new_G5214_ = ~new_G5210_;
  assign new_G1072_ = ~new_G5218_ | ~new_G5221_;
  assign new_G5222_ = ~new_G5218_;
  assign new_G1091_ = ~new_G5226_ | ~new_G5229_;
  assign new_G5230_ = ~new_G5226_;
  assign new_G1112_ = ~new_G1108_;
  assign new_G1121_ = ~new_G1117_;
  assign new_G1153_ = ~new_G5231_ | ~new_G5238_;
  assign new_G1157_ = ~new_G5239_ | ~new_G5246_;
  assign new_G5253_ = ~new_G5247_;
  assign new_G1216_ = ~new_G5247_ | ~new_G5254_;
  assign new_G5261_ = ~new_G5255_;
  assign new_G5262_ = ~new_G5258_;
  assign new_G5269_ = ~new_G5263_;
  assign new_G5270_ = ~new_G5266_;
  assign new_G5287_ = ~new_G5281_;
  assign new_G1239_ = ~new_G5281_ | ~new_G5288_;
  assign new_G5295_ = ~new_G5289_;
  assign new_G5296_ = ~new_G5292_;
  assign new_G5303_ = ~new_G5297_;
  assign new_G5304_ = ~new_G5300_;
  assign new_G5321_ = ~new_G5315_;
  assign new_G1262_ = ~new_G5315_ | ~new_G5322_;
  assign new_G5329_ = ~new_G5323_;
  assign new_G5330_ = ~new_G5326_;
  assign new_G5337_ = ~new_G5331_;
  assign new_G5338_ = ~new_G5334_;
  assign new_G1544_ = ~new_G5396_ | ~new_G5399_;
  assign new_G5400_ = ~new_G5396_;
  assign new_G1554_ = ~new_G5404_ | ~new_G5407_;
  assign new_G5408_ = ~new_G5404_;
  assign new_G1571_ = ~new_G5412_ | ~new_G5415_;
  assign new_G5416_ = ~new_G5412_;
  assign new_G1596_ = ~new_G5420_ | ~new_G5423_;
  assign new_G5424_ = ~new_G5420_;
  assign new_G1607_ = ~new_G5428_ | ~new_G5431_;
  assign new_G5432_ = ~new_G5428_;
  assign new_G1628_ = ~new_G5436_ | ~new_G5439_;
  assign new_G5440_ = ~new_G5436_;
  assign new_G1653_ = ~new_G5444_ | ~new_G5447_;
  assign new_G5448_ = ~new_G5444_;
  assign new_G1685_ = ~new_G5452_ | ~new_G5455_;
  assign new_G5456_ = ~new_G5452_;
  assign new_G1693_ = ~new_G5460_ | ~new_G5463_;
  assign new_G5464_ = ~new_G5460_;
  assign new_G1793_ = ~new_G5748_ | ~new_G5751_;
  assign new_G5752_ = ~new_G5748_;
  assign new_G1803_ = ~new_G5756_ | ~new_G5759_;
  assign new_G5760_ = ~new_G5756_;
  assign new_G1820_ = ~new_G5764_ | ~new_G5767_;
  assign new_G5768_ = ~new_G5764_;
  assign new_G1848_ = ~new_G5772_ | ~new_G5775_;
  assign new_G5776_ = ~new_G5772_;
  assign new_G1857_ = ~new_G5780_ | ~new_G5783_;
  assign new_G5784_ = ~new_G5780_;
  assign new_G1867_ = ~new_G5788_ | ~new_G5791_;
  assign new_G5792_ = ~new_G5788_;
  assign new_G1883_ = ~new_G5796_ | ~new_G5799_;
  assign new_G5800_ = ~new_G5796_;
  assign new_G1901_ = ~new_G5804_ | ~new_G5807_;
  assign new_G5808_ = ~new_G5804_;
  assign new_G1919_ = ~new_G5812_ | ~new_G5815_;
  assign new_G5816_ = ~new_G5812_;
  assign new_G5855_ = ~new_G5849_;
  assign new_G2351_ = new_G3751_ & new_G2111_;
  assign new_G2366_ = new_G3745_ & new_G2105_;
  assign new_G2384_ = new_G3739_ & new_G2099_;
  assign new_G2391_ = new_G2091_ & new_G3731_;
  assign new_G2417_ = new_G3725_ & new_G2085_;
  assign new_G2431_ = new_G3719_ & new_G2335_;
  assign new_G2448_ = new_G3713_ & new_G2329_;
  assign new_G2465_ = new_G3707_ & new_G2323_;
  assign new_G5935_ = ~new_G5929_;
  assign new_G2597_ = new_G3751_ & new_G2111_;
  assign new_G2612_ = new_G3745_ & new_G2105_;
  assign new_G2629_ = new_G3739_ & new_G2099_;
  assign new_G2635_ = new_G3731_ & new_G2091_;
  assign new_G2652_ = new_G3725_ & new_G2085_;
  assign new_G2670_ = new_G3719_ & new_G2335_;
  assign new_G2693_ = new_G3713_ & new_G2329_;
  assign new_G2715_ = new_G3707_ & new_G2323_;
  assign new_G6055_ = ~new_G6049_;
  assign new_G6373_ = ~new_G6367_;
  assign new_G6374_ = ~new_G6370_;
  assign new_G6381_ = ~new_G6375_;
  assign new_G6382_ = ~new_G6378_;
  assign new_G6389_ = ~new_G6383_;
  assign new_G6390_ = ~new_G6386_;
  assign new_G6397_ = ~new_G6391_;
  assign new_G6398_ = ~new_G6394_;
  assign new_G6405_ = ~new_G6399_;
  assign new_G6406_ = ~new_G6402_;
  assign new_G6413_ = ~new_G6407_;
  assign new_G6414_ = ~new_G6410_;
  assign new_G6421_ = ~new_G6415_;
  assign new_G6422_ = ~new_G6418_;
  assign new_G6429_ = ~new_G6423_;
  assign new_G6430_ = ~new_G6426_;
  assign new_G6437_ = ~new_G6431_;
  assign new_G6438_ = ~new_G6434_;
  assign new_G6446_ = ~new_G6442_;
  assign new_G3059_ = new_G4175_ & new_G3813_;
  assign new_G6454_ = ~new_G6450_;
  assign new_G3068_ = new_G4172_ & new_G3810_;
  assign new_G6462_ = ~new_G6458_;
  assign new_G3076_ = new_G4169_ & new_G3807_;
  assign new_G3079_ = new_G4166_ & new_G3804_;
  assign new_G6470_ = ~new_G6466_;
  assign new_G3090_ = new_G4163_ & new_G3801_;
  assign new_G3099_ = new_G4160_ & new_G2175_;
  assign new_G3107_ = new_G4157_ & new_G2171_;
  assign new_G3114_ = new_G4154_ & new_G2167_;
  assign new_G3116_ = new_G4151_ & new_G2163_;
  assign new_G6502_ = ~new_G6498_;
  assign new_G6525_ = ~new_G6519_;
  assign new_G6526_ = ~new_G6522_;
  assign new_G6533_ = ~new_G6527_;
  assign new_G6534_ = ~new_G6530_;
  assign new_G6541_ = ~new_G6535_;
  assign new_G6542_ = ~new_G6538_;
  assign new_G6549_ = ~new_G6543_;
  assign new_G6550_ = ~new_G6546_;
  assign new_G6565_ = ~new_G6559_;
  assign new_G6566_ = ~new_G6562_;
  assign new_G3220_ = ~new_G3216_;
  assign new_G3292_ = new_G4439_ & new_G3838_;
  assign new_G3308_ = new_G4434_ & new_G3833_;
  assign new_G3327_ = new_G4429_ & new_G3828_;
  assign new_G3335_ = new_G3821_ & new_G4422_;
  assign new_G3362_ = new_G4417_ & new_G3816_;
  assign new_G3376_ = new_G4412_ & new_G2198_;
  assign new_G3393_ = new_G4407_ & new_G2192_;
  assign new_G3410_ = new_G4402_ & new_G2186_;
  assign new_G3425_ = new_G4396_ & new_G2179_;
  assign new_G6693_ = ~new_G6687_;
  assign new_G3503_ = ~new_G6687_ | ~new_G6694_;
  assign new_G6701_ = ~new_G6695_;
  assign new_G6702_ = ~new_G6698_;
  assign new_G6709_ = ~new_G6703_;
  assign new_G6710_ = ~new_G6706_;
  assign new_G6728_ = ~new_G6724_;
  assign new_G6772_ = ~new_G6768_;
  assign new_G3853_ = new_G4439_ & new_G3838_;
  assign new_G3868_ = new_G4434_ & new_G3833_;
  assign new_G3885_ = new_G4429_ & new_G3828_;
  assign new_G3891_ = new_G4422_ & new_G3821_;
  assign new_G3908_ = new_G4417_ & new_G3816_;
  assign new_G3926_ = new_G4412_ & new_G2198_;
  assign new_G3949_ = new_G4407_ & new_G2192_;
  assign new_G3971_ = new_G4402_ & new_G2186_;
  assign new_G3979_ = new_G4396_ & new_G2179_;
  assign new_G7212_ = ~new_G7208_;
  assign new_G7227_ = ~new_G7221_;
  assign new_G7255_ = ~new_G7249_;
  assign new_G4202_ = ~new_G7249_ | ~new_G7256_;
  assign new_G7263_ = ~new_G7257_;
  assign new_G7264_ = ~new_G7260_;
  assign new_G7272_ = ~new_G7268_;
  assign new_G7299_ = ~new_G7293_;
  assign new_G4225_ = ~new_G7293_ | ~new_G7300_;
  assign new_G7307_ = ~new_G7301_;
  assign new_G7308_ = ~new_G7304_;
  assign new_G7315_ = ~new_G7309_;
  assign new_G7316_ = ~new_G7312_;
  assign new_G4297_ = new_G4511_ & new_G2081_;
  assign new_G4305_ = new_G4508_ & new_G2077_;
  assign new_G4312_ = new_G4505_ & new_G2073_;
  assign new_G4314_ = new_G4502_ & new_G2069_;
  assign new_G4324_ = new_G4499_ & new_G2065_;
  assign new_G7400_ = ~new_G7396_;
  assign new_G4333_ = new_G4496_ & new_G2316_;
  assign new_G7408_ = ~new_G7404_;
  assign new_G4341_ = new_G4493_ & new_G2312_;
  assign new_G7416_ = ~new_G7412_;
  assign new_G4348_ = new_G4490_ & new_G2308_;
  assign new_G4349_ = new_G3686_ & new_G3695_;
  assign new_G7431_ = ~new_G7425_;
  assign new_G4389_ = new_G2320_ & new_G1535_;
  assign new_G7469_ = ~new_G7463_;
  assign new_G4530_ = ~new_G7463_ | ~new_G7470_;
  assign new_G7477_ = ~new_G7471_;
  assign new_G7478_ = ~new_G7474_;
  assign new_G7485_ = ~new_G7479_;
  assign new_G7486_ = ~new_G7482_;
  assign new_G7513_ = ~new_G7507_;
  assign new_G7514_ = ~new_G7510_;
  assign new_G7558_ = ~new_G7554_;
  assign new_G4932_ = new_G917_ | new_G953_;
  assign new_G4956_ = ~new_G4952_;
  assign new_G4973_ = ~new_G917_;
  assign new_G4987_ = ~new_G4983_;
  assign new_G4997_ = ~new_G4993_;
  assign new_G5017_ = ~new_G5011_;
  assign new_G5099_ = new_G877_;
  assign new_G5345_ = ~new_G5339_;
  assign new_G5346_ = ~new_G5342_;
  assign new_G5355_ = ~new_G5349_;
  assign new_G5356_ = ~new_G5352_;
  assign new_G5372_ = ~new_G5279_ | ~new_G5280_;
  assign new_G5380_ = ~new_G5313_ | ~new_G5314_;
  assign new_G5471_ = ~new_G5465_;
  assign new_G5523_ = new_G1590_;
  assign new_G5587_ = ~new_G5581_;
  assign new_G5669_ = new_G1677_;
  assign new_G5857_ = new_G1841_;
  assign new_G5868_ = new_G2111_;
  assign new_G5876_ = new_G2105_;
  assign new_G5884_ = new_G2099_;
  assign new_G5892_ = new_G2091_;
  assign new_G5900_ = new_G2085_;
  assign new_G5908_ = new_G2335_;
  assign new_G5916_ = new_G2329_;
  assign new_G5924_ = new_G2323_;
  assign new_G5969_ = ~new_G2091_ & ~new_G3731_;
  assign new_G5988_ = new_G2111_;
  assign new_G5996_ = new_G2105_;
  assign new_G6004_ = new_G2099_;
  assign new_G6012_ = new_G2085_;
  assign new_G6020_ = new_G2335_;
  assign new_G6028_ = new_G2329_;
  assign new_G6036_ = new_G2323_;
  assign new_G6044_ = new_G2091_;
  assign new_G6057_ = ~new_G3731_ & ~new_G2091_;
  assign new_G6439_ = new_G4175_;
  assign new_G6447_ = new_G4172_;
  assign new_G6455_ = new_G4169_;
  assign new_G6463_ = new_G4163_;
  assign new_G6471_ = new_G4160_;
  assign new_G6474_ = new_G2175_;
  assign new_G6479_ = new_G4157_;
  assign new_G6482_ = new_G2171_;
  assign new_G6487_ = new_G4154_;
  assign new_G6490_ = new_G2167_;
  assign new_G6495_ = new_G4166_;
  assign new_G6503_ = new_G4151_;
  assign new_G6506_ = new_G2163_;
  assign new_G6570_ = new_G3838_;
  assign new_G6578_ = new_G3833_;
  assign new_G6586_ = new_G3828_;
  assign new_G6594_ = new_G3821_;
  assign new_G6602_ = new_G3816_;
  assign new_G6610_ = new_G2198_;
  assign new_G6618_ = new_G2192_;
  assign new_G6626_ = new_G2186_;
  assign new_G6634_ = new_G2179_;
  assign new_G6671_ = ~new_G3821_ & ~new_G4422_;
  assign new_G6721_ = new_G2179_;
  assign new_G6729_ = new_G2192_;
  assign new_G6732_ = new_G2186_;
  assign new_G6737_ = new_G3816_;
  assign new_G6740_ = new_G2198_;
  assign new_G6745_ = new_G3828_;
  assign new_G6748_ = new_G3821_;
  assign new_G6755_ = new_G3838_;
  assign new_G6758_ = new_G3833_;
  assign new_G6765_ = new_G2320_;
  assign new_G6773_ = new_G2329_;
  assign new_G6776_ = new_G2323_;
  assign new_G6781_ = new_G2085_;
  assign new_G6784_ = new_G2335_;
  assign new_G6789_ = new_G2099_;
  assign new_G6792_ = new_G2091_;
  assign new_G6799_ = new_G2111_;
  assign new_G6802_ = new_G2105_;
  assign new_G6832_ = ~new_G6719_ | ~new_G6720_;
  assign new_G6856_ = new_G3838_;
  assign new_G6864_ = new_G3833_;
  assign new_G6872_ = new_G3828_;
  assign new_G6880_ = new_G3816_;
  assign new_G6888_ = new_G2198_;
  assign new_G6896_ = new_G2192_;
  assign new_G6904_ = new_G2186_;
  assign new_G6912_ = new_G3821_;
  assign new_G6920_ = new_G2179_;
  assign new_G6925_ = ~new_G4422_ & ~new_G3821_;
  assign new_G7041_ = ~new_G4396_ & ~new_G2179_;
  assign new_G7205_ = new_G2163_;
  assign new_G7213_ = new_G2171_;
  assign new_G7216_ = new_G2167_;
  assign new_G7224_ = new_G2175_;
  assign new_G7235_ = ~new_G7229_;
  assign new_G7236_ = ~new_G7232_;
  assign new_G7245_ = ~new_G7239_;
  assign new_G7246_ = ~new_G7242_;
  assign new_G7265_ = new_G2065_;
  assign new_G7273_ = new_G2073_;
  assign new_G7276_ = new_G2069_;
  assign new_G7283_ = new_G2081_;
  assign new_G7286_ = new_G2077_;
  assign new_G7323_ = ~new_G7317_;
  assign new_G7324_ = ~new_G7320_;
  assign new_G7333_ = ~new_G7327_;
  assign new_G7334_ = ~new_G7330_;
  assign new_G7361_ = new_G4511_;
  assign new_G7364_ = new_G2081_;
  assign new_G7369_ = new_G4508_;
  assign new_G7372_ = new_G2077_;
  assign new_G7377_ = new_G4505_;
  assign new_G7380_ = new_G2073_;
  assign new_G7385_ = new_G4499_;
  assign new_G7388_ = new_G2065_;
  assign new_G7393_ = new_G4496_;
  assign new_G7401_ = new_G4493_;
  assign new_G7409_ = new_G4490_;
  assign new_G7417_ = new_G4502_;
  assign new_G7420_ = new_G2069_;
  assign new_G7428_ = new_G3695_;
  assign new_G7493_ = ~new_G7487_;
  assign new_G7494_ = ~new_G7490_;
  assign new_G7503_ = ~new_G7497_;
  assign new_G7504_ = ~new_G7500_;
  assign new_G7515_ = new_G4493_;
  assign new_G7518_ = new_G4490_;
  assign new_G7523_ = new_G4499_;
  assign new_G7526_ = new_G4496_;
  assign new_G7531_ = new_G4505_;
  assign new_G7534_ = new_G4502_;
  assign new_G7541_ = new_G4511_;
  assign new_G7544_ = new_G4508_;
  assign new_G7551_ = new_G4151_;
  assign new_G7559_ = new_G4157_;
  assign new_G7562_ = new_G4154_;
  assign new_G7567_ = new_G4163_;
  assign new_G7570_ = new_G4160_;
  assign new_G7575_ = new_G4169_;
  assign new_G7578_ = new_G4166_;
  assign new_G7585_ = new_G4175_;
  assign new_G7588_ = new_G4172_;
  assign new_G1176_ = ~new_G1121_ | ~new_G1112_;
  assign new_G957_ = ~new_G912_ | ~new_G906_;
  assign new_G791_ = ~new_G4881_ | ~new_G4888_;
  assign new_G804_ = ~new_G4889_ | ~new_G4896_;
  assign new_G826_ = ~new_G4897_ | ~new_G4904_;
  assign new_G852_ = ~new_G4905_ | ~new_G4912_;
  assign new_G894_ = ~new_G4921_ | ~new_G4928_;
  assign new_G1025_ = ~new_G5191_ | ~new_G5198_;
  assign new_G1037_ = ~new_G5199_ | ~new_G5206_;
  assign new_G1054_ = ~new_G5207_ | ~new_G5214_;
  assign new_G1073_ = ~new_G5215_ | ~new_G5222_;
  assign new_G1092_ = ~new_G5223_ | ~new_G5230_;
  assign new_G1154_ = ~new_G1152_ | ~new_G1153_;
  assign new_G1158_ = ~new_G1156_ | ~new_G1157_;
  assign new_G1215_ = ~new_G5250_ | ~new_G5253_;
  assign new_G1224_ = ~new_G5258_ | ~new_G5261_;
  assign new_G1225_ = ~new_G5255_ | ~new_G5262_;
  assign new_G1233_ = ~new_G5266_ | ~new_G5269_;
  assign new_G1234_ = ~new_G5263_ | ~new_G5270_;
  assign new_G1238_ = ~new_G5284_ | ~new_G5287_;
  assign new_G1247_ = ~new_G5292_ | ~new_G5295_;
  assign new_G1248_ = ~new_G5289_ | ~new_G5296_;
  assign new_G1256_ = ~new_G5300_ | ~new_G5303_;
  assign new_G1257_ = ~new_G5297_ | ~new_G5304_;
  assign new_G1261_ = ~new_G5318_ | ~new_G5321_;
  assign new_G1270_ = ~new_G5326_ | ~new_G5329_;
  assign new_G1271_ = ~new_G5323_ | ~new_G5330_;
  assign new_G1279_ = ~new_G5334_ | ~new_G5337_;
  assign new_G1280_ = ~new_G5331_ | ~new_G5338_;
  assign new_G1545_ = ~new_G5393_ | ~new_G5400_;
  assign new_G1555_ = ~new_G5401_ | ~new_G5408_;
  assign new_G1572_ = ~new_G5409_ | ~new_G5416_;
  assign new_G1597_ = ~new_G5417_ | ~new_G5424_;
  assign new_G1608_ = ~new_G5425_ | ~new_G5432_;
  assign new_G1629_ = ~new_G5433_ | ~new_G5440_;
  assign new_G1654_ = ~new_G5441_ | ~new_G5448_;
  assign new_G1686_ = ~new_G5449_ | ~new_G5456_;
  assign new_G1694_ = ~new_G5457_ | ~new_G5464_;
  assign new_G1794_ = ~new_G5745_ | ~new_G5752_;
  assign new_G1804_ = ~new_G5753_ | ~new_G5760_;
  assign new_G1821_ = ~new_G5761_ | ~new_G5768_;
  assign new_G1849_ = ~new_G5769_ | ~new_G5776_;
  assign new_G1858_ = ~new_G5777_ | ~new_G5784_;
  assign new_G1868_ = ~new_G5785_ | ~new_G5792_;
  assign new_G1884_ = ~new_G5793_ | ~new_G5800_;
  assign new_G1902_ = ~new_G5801_ | ~new_G5808_;
  assign new_G1920_ = ~new_G5809_ | ~new_G5816_;
  assign new_G2954_ = ~new_G6370_ | ~new_G6373_;
  assign new_G2955_ = ~new_G6367_ | ~new_G6374_;
  assign new_G2963_ = ~new_G6378_ | ~new_G6381_;
  assign new_G2964_ = ~new_G6375_ | ~new_G6382_;
  assign new_G2971_ = ~new_G6386_ | ~new_G6389_;
  assign new_G2972_ = ~new_G6383_ | ~new_G6390_;
  assign new_G2980_ = ~new_G6394_ | ~new_G6397_;
  assign new_G2981_ = ~new_G6391_ | ~new_G6398_;
  assign new_G2990_ = ~new_G6402_ | ~new_G6405_;
  assign new_G2991_ = ~new_G6399_ | ~new_G6406_;
  assign new_G2999_ = ~new_G6410_ | ~new_G6413_;
  assign new_G3000_ = ~new_G6407_ | ~new_G6414_;
  assign new_G3007_ = ~new_G6418_ | ~new_G6421_;
  assign new_G3008_ = ~new_G6415_ | ~new_G6422_;
  assign new_G3016_ = ~new_G6426_ | ~new_G6429_;
  assign new_G3017_ = ~new_G6423_ | ~new_G6430_;
  assign new_G3019_ = ~new_G6434_ | ~new_G6437_;
  assign new_G3020_ = ~new_G6431_ | ~new_G6438_;
  assign new_G3174_ = ~new_G6522_ | ~new_G6525_;
  assign new_G3175_ = ~new_G6519_ | ~new_G6526_;
  assign new_G3184_ = ~new_G6530_ | ~new_G6533_;
  assign new_G3185_ = ~new_G6527_ | ~new_G6534_;
  assign new_G3193_ = ~new_G6538_ | ~new_G6541_;
  assign new_G3194_ = ~new_G6535_ | ~new_G6542_;
  assign new_G3201_ = ~new_G6546_ | ~new_G6549_;
  assign new_G3202_ = ~new_G6543_ | ~new_G6550_;
  assign new_G3213_ = ~new_G6562_ | ~new_G6565_;
  assign new_G3214_ = ~new_G6559_ | ~new_G6566_;
  assign new_G3227_ = ~new_G3223_;
  assign new_G3502_ = ~new_G6690_ | ~new_G6693_;
  assign new_G3511_ = ~new_G6698_ | ~new_G6701_;
  assign new_G3512_ = ~new_G6695_ | ~new_G6702_;
  assign new_G3520_ = ~new_G6706_ | ~new_G6709_;
  assign new_G3521_ = ~new_G6703_ | ~new_G6710_;
  assign new_G4201_ = ~new_G7252_ | ~new_G7255_;
  assign new_G4210_ = ~new_G7260_ | ~new_G7263_;
  assign new_G4211_ = ~new_G7257_ | ~new_G7264_;
  assign new_G4224_ = ~new_G7296_ | ~new_G7299_;
  assign new_G4233_ = ~new_G7304_ | ~new_G7307_;
  assign new_G4234_ = ~new_G7301_ | ~new_G7308_;
  assign new_G4242_ = ~new_G7312_ | ~new_G7315_;
  assign new_G4243_ = ~new_G7309_ | ~new_G7316_;
  assign new_G4529_ = ~new_G7466_ | ~new_G7469_;
  assign new_G4538_ = ~new_G7474_ | ~new_G7477_;
  assign new_G4539_ = ~new_G7471_ | ~new_G7478_;
  assign new_G4547_ = ~new_G7482_ | ~new_G7485_;
  assign new_G4548_ = ~new_G7479_ | ~new_G7486_;
  assign new_G4552_ = ~new_G7510_ | ~new_G7513_;
  assign new_G4553_ = ~new_G7507_ | ~new_G7514_;
  assign new_G4946_ = ~new_G4942_;
  assign new_G5347_ = ~new_G5342_ | ~new_G5345_;
  assign new_G5348_ = ~new_G5339_ | ~new_G5346_;
  assign new_G5357_ = ~new_G5352_ | ~new_G5355_;
  assign new_G5358_ = ~new_G5349_ | ~new_G5356_;
  assign new_G7237_ = ~new_G7232_ | ~new_G7235_;
  assign new_G7238_ = ~new_G7229_ | ~new_G7236_;
  assign new_G7247_ = ~new_G7242_ | ~new_G7245_;
  assign new_G7248_ = ~new_G7239_ | ~new_G7246_;
  assign new_G7325_ = ~new_G7320_ | ~new_G7323_;
  assign new_G7326_ = ~new_G7317_ | ~new_G7324_;
  assign new_G7335_ = ~new_G7330_ | ~new_G7333_;
  assign new_G7336_ = ~new_G7327_ | ~new_G7334_;
  assign new_G7495_ = ~new_G7490_ | ~new_G7493_;
  assign new_G7496_ = ~new_G7487_ | ~new_G7494_;
  assign new_G7505_ = ~new_G7500_ | ~new_G7503_;
  assign new_G7506_ = ~new_G7497_ | ~new_G7504_;
  assign new_G3244_ = ~new_G3227_ | ~new_G3220_;
  assign new_G792_ = ~new_G790_ | ~new_G791_;
  assign new_G805_ = ~new_G803_ | ~new_G804_;
  assign new_G827_ = ~new_G825_ | ~new_G826_;
  assign new_G853_ = ~new_G851_ | ~new_G852_;
  assign new_G895_ = ~new_G893_ | ~new_G894_;
  assign new_G1026_ = ~new_G1024_ | ~new_G1025_;
  assign new_G1038_ = ~new_G1036_ | ~new_G1037_;
  assign new_G1055_ = ~new_G1053_ | ~new_G1054_;
  assign new_G1074_ = ~new_G1072_ | ~new_G1073_;
  assign new_G1093_ = ~new_G1091_ | ~new_G1092_;
  assign new_G1155_ = ~new_G1154_;
  assign new_G1217_ = ~new_G1215_ | ~new_G1216_;
  assign new_G1226_ = ~new_G1224_ | ~new_G1225_;
  assign new_G1235_ = ~new_G1233_ | ~new_G1234_;
  assign new_G1240_ = ~new_G1238_ | ~new_G1239_;
  assign new_G1249_ = ~new_G1247_ | ~new_G1248_;
  assign new_G1258_ = ~new_G1256_ | ~new_G1257_;
  assign new_G1263_ = ~new_G1261_ | ~new_G1262_;
  assign new_G1272_ = ~new_G1270_ | ~new_G1271_;
  assign new_G1281_ = ~new_G1279_ | ~new_G1280_;
  assign new_G5376_ = ~new_G5372_;
  assign new_G5384_ = ~new_G5380_;
  assign new_G1546_ = ~new_G1544_ | ~new_G1545_;
  assign new_G1556_ = ~new_G1554_ | ~new_G1555_;
  assign new_G1573_ = ~new_G1571_ | ~new_G1572_;
  assign new_G1598_ = ~new_G1596_ | ~new_G1597_;
  assign new_G1609_ = ~new_G1607_ | ~new_G1608_;
  assign new_G1630_ = ~new_G1628_ | ~new_G1629_;
  assign new_G1655_ = ~new_G1653_ | ~new_G1654_;
  assign new_G1687_ = ~new_G1685_ | ~new_G1686_;
  assign new_G1695_ = ~new_G1693_ | ~new_G1694_;
  assign new_G1795_ = ~new_G1793_ | ~new_G1794_;
  assign new_G1805_ = ~new_G1803_ | ~new_G1804_;
  assign new_G1822_ = ~new_G1820_ | ~new_G1821_;
  assign new_G1850_ = ~new_G1848_ | ~new_G1849_;
  assign new_G1859_ = ~new_G1857_ | ~new_G1858_;
  assign new_G1869_ = ~new_G1867_ | ~new_G1868_;
  assign new_G1885_ = ~new_G1883_ | ~new_G1884_;
  assign new_G1903_ = ~new_G1901_ | ~new_G1902_;
  assign new_G1921_ = ~new_G1919_ | ~new_G1920_;
  assign new_G5863_ = ~new_G5857_;
  assign new_G2341_ = ~new_G5868_ | ~new_G5871_;
  assign new_G5872_ = ~new_G5868_;
  assign new_G2352_ = ~new_G5876_ | ~new_G5879_;
  assign new_G5880_ = ~new_G5876_;
  assign new_G2370_ = ~new_G5884_ | ~new_G5887_;
  assign new_G5888_ = ~new_G5884_;
  assign new_G2398_ = ~new_G5892_ | ~new_G5895_;
  assign new_G5896_ = ~new_G5892_;
  assign new_G2407_ = ~new_G5900_ | ~new_G5903_;
  assign new_G5904_ = ~new_G5900_;
  assign new_G2418_ = ~new_G5908_ | ~new_G5911_;
  assign new_G5912_ = ~new_G5908_;
  assign new_G2434_ = ~new_G5916_ | ~new_G5919_;
  assign new_G5920_ = ~new_G5916_;
  assign new_G2452_ = ~new_G5924_ | ~new_G5927_;
  assign new_G5928_ = ~new_G5924_;
  assign new_G2481_ = new_G3682_ & new_G4389_;
  assign new_G5975_ = ~new_G5969_;
  assign new_G2587_ = ~new_G5988_ | ~new_G5991_;
  assign new_G5992_ = ~new_G5988_;
  assign new_G2598_ = ~new_G5996_ | ~new_G5999_;
  assign new_G6000_ = ~new_G5996_;
  assign new_G2616_ = ~new_G6004_ | ~new_G6007_;
  assign new_G6008_ = ~new_G6004_;
  assign new_G2641_ = ~new_G6012_ | ~new_G6015_;
  assign new_G6016_ = ~new_G6012_;
  assign new_G2653_ = ~new_G6020_ | ~new_G6023_;
  assign new_G6024_ = ~new_G6020_;
  assign new_G2674_ = ~new_G6028_ | ~new_G6031_;
  assign new_G6032_ = ~new_G6028_;
  assign new_G2699_ = ~new_G6036_ | ~new_G6039_;
  assign new_G6040_ = ~new_G6036_;
  assign new_G2724_ = new_G3682_ & new_G4389_;
  assign new_G2732_ = ~new_G6044_ | ~new_G6047_;
  assign new_G6048_ = ~new_G6044_;
  assign new_G2956_ = ~new_G2954_ | ~new_G2955_;
  assign new_G2965_ = ~new_G2963_ | ~new_G2964_;
  assign new_G2973_ = ~new_G2971_ | ~new_G2972_;
  assign new_G2982_ = ~new_G2980_ | ~new_G2981_;
  assign new_G2992_ = ~new_G2990_ | ~new_G2991_;
  assign new_G3001_ = ~new_G2999_ | ~new_G3000_;
  assign new_G3009_ = ~new_G3007_ | ~new_G3008_;
  assign new_G3018_ = ~new_G3016_ | ~new_G3017_;
  assign new_G3021_ = ~new_G3019_ | ~new_G3020_;
  assign new_G6445_ = ~new_G6439_;
  assign new_G3051_ = ~new_G6439_ | ~new_G6446_;
  assign new_G6453_ = ~new_G6447_;
  assign new_G3061_ = ~new_G6447_ | ~new_G6454_;
  assign new_G6461_ = ~new_G6455_;
  assign new_G3070_ = ~new_G6455_ | ~new_G6462_;
  assign new_G6469_ = ~new_G6463_;
  assign new_G3081_ = ~new_G6463_ | ~new_G6470_;
  assign new_G6477_ = ~new_G6471_;
  assign new_G6478_ = ~new_G6474_;
  assign new_G6485_ = ~new_G6479_;
  assign new_G6486_ = ~new_G6482_;
  assign new_G6493_ = ~new_G6487_;
  assign new_G6494_ = ~new_G6490_;
  assign new_G6501_ = ~new_G6495_;
  assign new_G3118_ = ~new_G6495_ | ~new_G6502_;
  assign new_G6509_ = ~new_G6503_;
  assign new_G6510_ = ~new_G6506_;
  assign new_G3176_ = ~new_G3174_ | ~new_G3175_;
  assign new_G3186_ = ~new_G3184_ | ~new_G3185_;
  assign new_G3195_ = ~new_G3193_ | ~new_G3194_;
  assign new_G3203_ = ~new_G3201_ | ~new_G3202_;
  assign new_G3215_ = ~new_G3213_ | ~new_G3214_;
  assign new_G3281_ = ~new_G6570_ | ~new_G6573_;
  assign new_G6574_ = ~new_G6570_;
  assign new_G3293_ = ~new_G6578_ | ~new_G6581_;
  assign new_G6582_ = ~new_G6578_;
  assign new_G3312_ = ~new_G6586_ | ~new_G6589_;
  assign new_G6590_ = ~new_G6586_;
  assign new_G3342_ = ~new_G6594_ | ~new_G6597_;
  assign new_G6598_ = ~new_G6594_;
  assign new_G3351_ = ~new_G6602_ | ~new_G6605_;
  assign new_G6606_ = ~new_G6602_;
  assign new_G3363_ = ~new_G6610_ | ~new_G6613_;
  assign new_G6614_ = ~new_G6610_;
  assign new_G3379_ = ~new_G6618_ | ~new_G6621_;
  assign new_G6622_ = ~new_G6618_;
  assign new_G3397_ = ~new_G6626_ | ~new_G6629_;
  assign new_G6630_ = ~new_G6626_;
  assign new_G3415_ = ~new_G6634_ | ~new_G6637_;
  assign new_G6638_ = ~new_G6634_;
  assign new_G6677_ = ~new_G6671_;
  assign new_G3504_ = ~new_G3502_ | ~new_G3503_;
  assign new_G3513_ = ~new_G3511_ | ~new_G3512_;
  assign new_G3522_ = ~new_G3520_ | ~new_G3521_;
  assign new_G6727_ = ~new_G6721_;
  assign new_G3526_ = ~new_G6721_ | ~new_G6728_;
  assign new_G6735_ = ~new_G6729_;
  assign new_G6736_ = ~new_G6732_;
  assign new_G6743_ = ~new_G6737_;
  assign new_G6744_ = ~new_G6740_;
  assign new_G6771_ = ~new_G6765_;
  assign new_G3549_ = ~new_G6765_ | ~new_G6772_;
  assign new_G6779_ = ~new_G6773_;
  assign new_G6780_ = ~new_G6776_;
  assign new_G6787_ = ~new_G6781_;
  assign new_G6788_ = ~new_G6784_;
  assign new_G6836_ = ~new_G6832_;
  assign new_G3843_ = ~new_G6856_ | ~new_G6859_;
  assign new_G6860_ = ~new_G6856_;
  assign new_G3854_ = ~new_G6864_ | ~new_G6867_;
  assign new_G6868_ = ~new_G6864_;
  assign new_G3872_ = ~new_G6872_ | ~new_G6875_;
  assign new_G6876_ = ~new_G6872_;
  assign new_G3897_ = ~new_G6880_ | ~new_G6883_;
  assign new_G6884_ = ~new_G6880_;
  assign new_G3909_ = ~new_G6888_ | ~new_G6891_;
  assign new_G6892_ = ~new_G6888_;
  assign new_G3930_ = ~new_G6896_ | ~new_G6899_;
  assign new_G6900_ = ~new_G6896_;
  assign new_G3955_ = ~new_G6904_ | ~new_G6907_;
  assign new_G6908_ = ~new_G6904_;
  assign new_G3987_ = ~new_G6912_ | ~new_G6915_;
  assign new_G6916_ = ~new_G6912_;
  assign new_G3995_ = ~new_G6920_ | ~new_G6923_;
  assign new_G6924_ = ~new_G6920_;
  assign new_G7211_ = ~new_G7205_;
  assign new_G4179_ = ~new_G7205_ | ~new_G7212_;
  assign new_G7219_ = ~new_G7213_;
  assign new_G7220_ = ~new_G7216_;
  assign new_G4196_ = ~new_G7224_ | ~new_G7227_;
  assign new_G7228_ = ~new_G7224_;
  assign new_G4203_ = ~new_G4201_ | ~new_G4202_;
  assign new_G4212_ = ~new_G4210_ | ~new_G4211_;
  assign new_G7271_ = ~new_G7265_;
  assign new_G4220_ = ~new_G7265_ | ~new_G7272_;
  assign new_G4226_ = ~new_G4224_ | ~new_G4225_;
  assign new_G4235_ = ~new_G4233_ | ~new_G4234_;
  assign new_G4244_ = ~new_G4242_ | ~new_G4243_;
  assign new_G7367_ = ~new_G7361_;
  assign new_G7368_ = ~new_G7364_;
  assign new_G7375_ = ~new_G7369_;
  assign new_G7376_ = ~new_G7372_;
  assign new_G7383_ = ~new_G7377_;
  assign new_G7384_ = ~new_G7380_;
  assign new_G7391_ = ~new_G7385_;
  assign new_G7392_ = ~new_G7388_;
  assign new_G7399_ = ~new_G7393_;
  assign new_G4326_ = ~new_G7393_ | ~new_G7400_;
  assign new_G7407_ = ~new_G7401_;
  assign new_G4335_ = ~new_G7401_ | ~new_G7408_;
  assign new_G7415_ = ~new_G7409_;
  assign new_G4343_ = ~new_G7409_ | ~new_G7416_;
  assign new_G7423_ = ~new_G7417_;
  assign new_G7424_ = ~new_G7420_;
  assign new_G4353_ = ~new_G7428_ | ~new_G7431_;
  assign new_G7432_ = ~new_G7428_;
  assign new_G4531_ = ~new_G4529_ | ~new_G4530_;
  assign new_G4540_ = ~new_G4538_ | ~new_G4539_;
  assign new_G4549_ = ~new_G4547_ | ~new_G4548_;
  assign new_G4554_ = ~new_G4552_ | ~new_G4553_;
  assign new_G7521_ = ~new_G7515_;
  assign new_G7522_ = ~new_G7518_;
  assign new_G7529_ = ~new_G7523_;
  assign new_G7530_ = ~new_G7526_;
  assign new_G7557_ = ~new_G7551_;
  assign new_G4576_ = ~new_G7551_ | ~new_G7558_;
  assign new_G7565_ = ~new_G7559_;
  assign new_G7566_ = ~new_G7562_;
  assign new_G7573_ = ~new_G7567_;
  assign new_G7574_ = ~new_G7570_;
  assign new_G4936_ = ~new_G4932_;
  assign new_G4937_ = ~new_G4932_ | ~new_G4935_;
  assign new_G4977_ = ~new_G4973_;
  assign new_G4978_ = ~new_G4973_ | ~new_G4976_;
  assign new_G5105_ = ~new_G5099_;
  assign new_G5359_ = ~new_G5357_ | ~new_G5358_;
  assign new_G5362_ = ~new_G5347_ | ~new_G5348_;
  assign new_G5529_ = ~new_G5523_;
  assign new_G5675_ = ~new_G5669_;
  assign new_G5932_ = new_G4389_;
  assign new_G5977_ = new_G2391_;
  assign new_G6052_ = new_G4389_;
  assign new_G6063_ = ~new_G6057_;
  assign new_G6115_ = new_G2635_;
  assign new_G6173_ = ~new_G3682_ & ~new_G4389_;
  assign new_G6679_ = new_G3335_;
  assign new_G6751_ = ~new_G6745_;
  assign new_G6752_ = ~new_G6748_;
  assign new_G6761_ = ~new_G6755_;
  assign new_G6762_ = ~new_G6758_;
  assign new_G6795_ = ~new_G6789_;
  assign new_G6796_ = ~new_G6792_;
  assign new_G6805_ = ~new_G6799_;
  assign new_G6806_ = ~new_G6802_;
  assign new_G6931_ = ~new_G6925_;
  assign new_G6983_ = new_G3891_;
  assign new_G7047_ = ~new_G7041_;
  assign new_G7129_ = new_G3979_;
  assign new_G7279_ = ~new_G7273_;
  assign new_G7280_ = ~new_G7276_;
  assign new_G7289_ = ~new_G7283_;
  assign new_G7290_ = ~new_G7286_;
  assign new_G7337_ = ~new_G7247_ | ~new_G7248_;
  assign new_G7340_ = ~new_G7237_ | ~new_G7238_;
  assign new_G7353_ = ~new_G7335_ | ~new_G7336_;
  assign new_G7356_ = ~new_G7325_ | ~new_G7326_;
  assign new_G7537_ = ~new_G7531_;
  assign new_G7538_ = ~new_G7534_;
  assign new_G7547_ = ~new_G7541_;
  assign new_G7548_ = ~new_G7544_;
  assign new_G7581_ = ~new_G7575_;
  assign new_G7582_ = ~new_G7578_;
  assign new_G7591_ = ~new_G7585_;
  assign new_G7592_ = ~new_G7588_;
  assign new_G7595_ = ~new_G7505_ | ~new_G7506_;
  assign new_G7598_ = ~new_G7495_ | ~new_G7496_;
  assign new_G2342_ = ~new_G5865_ | ~new_G5872_;
  assign new_G2353_ = ~new_G5873_ | ~new_G5880_;
  assign new_G2371_ = ~new_G5881_ | ~new_G5888_;
  assign new_G2399_ = ~new_G5889_ | ~new_G5896_;
  assign new_G2408_ = ~new_G5897_ | ~new_G5904_;
  assign new_G2419_ = ~new_G5905_ | ~new_G5912_;
  assign new_G2435_ = ~new_G5913_ | ~new_G5920_;
  assign new_G2453_ = ~new_G5921_ | ~new_G5928_;
  assign new_G2588_ = ~new_G5985_ | ~new_G5992_;
  assign new_G2599_ = ~new_G5993_ | ~new_G6000_;
  assign new_G2617_ = ~new_G6001_ | ~new_G6008_;
  assign new_G2642_ = ~new_G6009_ | ~new_G6016_;
  assign new_G2654_ = ~new_G6017_ | ~new_G6024_;
  assign new_G2675_ = ~new_G6025_ | ~new_G6032_;
  assign new_G2700_ = ~new_G6033_ | ~new_G6040_;
  assign new_G2733_ = ~new_G6041_ | ~new_G6048_;
  assign new_G3050_ = ~new_G6442_ | ~new_G6445_;
  assign new_G3060_ = ~new_G6450_ | ~new_G6453_;
  assign new_G3069_ = ~new_G6458_ | ~new_G6461_;
  assign new_G3080_ = ~new_G6466_ | ~new_G6469_;
  assign new_G3091_ = ~new_G6474_ | ~new_G6477_;
  assign new_G3092_ = ~new_G6471_ | ~new_G6478_;
  assign new_G3100_ = ~new_G6482_ | ~new_G6485_;
  assign new_G3101_ = ~new_G6479_ | ~new_G6486_;
  assign new_G3108_ = ~new_G6490_ | ~new_G6493_;
  assign new_G3109_ = ~new_G6487_ | ~new_G6494_;
  assign new_G3117_ = ~new_G6498_ | ~new_G6501_;
  assign new_G3120_ = ~new_G6506_ | ~new_G6509_;
  assign new_G3121_ = ~new_G6503_ | ~new_G6510_;
  assign new_G3282_ = ~new_G6567_ | ~new_G6574_;
  assign new_G3294_ = ~new_G6575_ | ~new_G6582_;
  assign new_G3313_ = ~new_G6583_ | ~new_G6590_;
  assign new_G3343_ = ~new_G6591_ | ~new_G6598_;
  assign new_G3352_ = ~new_G6599_ | ~new_G6606_;
  assign new_G3364_ = ~new_G6607_ | ~new_G6614_;
  assign new_G3380_ = ~new_G6615_ | ~new_G6622_;
  assign new_G3398_ = ~new_G6623_ | ~new_G6630_;
  assign new_G3416_ = ~new_G6631_ | ~new_G6638_;
  assign new_G3525_ = ~new_G6724_ | ~new_G6727_;
  assign new_G3534_ = ~new_G6732_ | ~new_G6735_;
  assign new_G3535_ = ~new_G6729_ | ~new_G6736_;
  assign new_G3543_ = ~new_G6740_ | ~new_G6743_;
  assign new_G3544_ = ~new_G6737_ | ~new_G6744_;
  assign new_G3548_ = ~new_G6768_ | ~new_G6771_;
  assign new_G3557_ = ~new_G6776_ | ~new_G6779_;
  assign new_G3558_ = ~new_G6773_ | ~new_G6780_;
  assign new_G3566_ = ~new_G6784_ | ~new_G6787_;
  assign new_G3567_ = ~new_G6781_ | ~new_G6788_;
  assign new_G3844_ = ~new_G6853_ | ~new_G6860_;
  assign new_G3855_ = ~new_G6861_ | ~new_G6868_;
  assign new_G3873_ = ~new_G6869_ | ~new_G6876_;
  assign new_G3898_ = ~new_G6877_ | ~new_G6884_;
  assign new_G3910_ = ~new_G6885_ | ~new_G6892_;
  assign new_G3931_ = ~new_G6893_ | ~new_G6900_;
  assign new_G3956_ = ~new_G6901_ | ~new_G6908_;
  assign new_G3988_ = ~new_G6909_ | ~new_G6916_;
  assign new_G3996_ = ~new_G6917_ | ~new_G6924_;
  assign new_G4178_ = ~new_G7208_ | ~new_G7211_;
  assign new_G4187_ = ~new_G7216_ | ~new_G7219_;
  assign new_G4188_ = ~new_G7213_ | ~new_G7220_;
  assign new_G4197_ = ~new_G7221_ | ~new_G7228_;
  assign new_G4219_ = ~new_G7268_ | ~new_G7271_;
  assign new_G4289_ = ~new_G7364_ | ~new_G7367_;
  assign new_G4290_ = ~new_G7361_ | ~new_G7368_;
  assign new_G4298_ = ~new_G7372_ | ~new_G7375_;
  assign new_G4299_ = ~new_G7369_ | ~new_G7376_;
  assign new_G4306_ = ~new_G7380_ | ~new_G7383_;
  assign new_G4307_ = ~new_G7377_ | ~new_G7384_;
  assign new_G4315_ = ~new_G7388_ | ~new_G7391_;
  assign new_G4316_ = ~new_G7385_ | ~new_G7392_;
  assign new_G4325_ = ~new_G7396_ | ~new_G7399_;
  assign new_G4334_ = ~new_G7404_ | ~new_G7407_;
  assign new_G4342_ = ~new_G7412_ | ~new_G7415_;
  assign new_G4350_ = ~new_G7420_ | ~new_G7423_;
  assign new_G4351_ = ~new_G7417_ | ~new_G7424_;
  assign new_G4354_ = ~new_G7425_ | ~new_G7432_;
  assign new_G4561_ = ~new_G7518_ | ~new_G7521_;
  assign new_G4562_ = ~new_G7515_ | ~new_G7522_;
  assign new_G4570_ = ~new_G7526_ | ~new_G7529_;
  assign new_G4571_ = ~new_G7523_ | ~new_G7530_;
  assign new_G4575_ = ~new_G7554_ | ~new_G7557_;
  assign new_G4584_ = ~new_G7562_ | ~new_G7565_;
  assign new_G4585_ = ~new_G7559_ | ~new_G7566_;
  assign new_G4593_ = ~new_G7570_ | ~new_G7573_;
  assign new_G4594_ = ~new_G7567_ | ~new_G7574_;
  assign new_G4938_ = ~new_G4929_ | ~new_G4936_;
  assign new_G4979_ = ~new_G4970_ | ~new_G4977_;
  assign new_G6753_ = ~new_G6748_ | ~new_G6751_;
  assign new_G6754_ = ~new_G6745_ | ~new_G6752_;
  assign new_G6763_ = ~new_G6758_ | ~new_G6761_;
  assign new_G6764_ = ~new_G6755_ | ~new_G6762_;
  assign new_G6797_ = ~new_G6792_ | ~new_G6795_;
  assign new_G6798_ = ~new_G6789_ | ~new_G6796_;
  assign new_G6807_ = ~new_G6802_ | ~new_G6805_;
  assign new_G6808_ = ~new_G6799_ | ~new_G6806_;
  assign new_G7281_ = ~new_G7276_ | ~new_G7279_;
  assign new_G7282_ = ~new_G7273_ | ~new_G7280_;
  assign new_G7291_ = ~new_G7286_ | ~new_G7289_;
  assign new_G7292_ = ~new_G7283_ | ~new_G7290_;
  assign new_G7539_ = ~new_G7534_ | ~new_G7537_;
  assign new_G7540_ = ~new_G7531_ | ~new_G7538_;
  assign new_G7549_ = ~new_G7544_ | ~new_G7547_;
  assign new_G7550_ = ~new_G7541_ | ~new_G7548_;
  assign new_G7583_ = ~new_G7578_ | ~new_G7581_;
  assign new_G7584_ = ~new_G7575_ | ~new_G7582_;
  assign new_G7593_ = ~new_G7588_ | ~new_G7591_;
  assign new_G7594_ = ~new_G7585_ | ~new_G7592_;
  assign new_G1856_ = ~new_G1850_;
  assign new_G920_ = new_G792_ & new_G805_ & new_G827_ & new_G895_ & new_G853_;
  assign new_G925_ = new_G792_ & new_G821_;
  assign new_G926_ = new_G845_ & new_G805_ & new_G792_;
  assign new_G927_ = new_G805_ & new_G868_ & new_G827_ & new_G792_;
  assign new_G928_ = new_G805_ & new_G877_ & new_G792_ & new_G853_ & new_G827_;
  assign new_G937_ = new_G805_ & new_G845_;
  assign new_G938_ = new_G805_ & new_G827_ & new_G868_;
  assign new_G939_ = new_G805_ & new_G877_ & new_G853_ & new_G827_;
  assign new_G940_ = new_G853_ & new_G805_ & new_G895_ & new_G827_;
  assign new_G941_ = new_G805_ & new_G845_;
  assign new_G942_ = new_G805_ & new_G827_ & new_G868_;
  assign new_G943_ = new_G805_ & new_G877_ & new_G853_ & new_G827_;
  assign new_G944_ = new_G827_ & new_G868_;
  assign new_G945_ = new_G877_ & new_G853_ & new_G827_;
  assign new_G946_ = new_G853_ & new_G895_ & new_G827_;
  assign new_G947_ = new_G827_ & new_G868_;
  assign new_G948_ = new_G877_ & new_G853_ & new_G827_;
  assign new_G949_ = new_G853_ & new_G877_;
  assign new_G956_ = new_G895_ & new_G853_;
  assign new_G1122_ = new_G1074_ & new_G1026_ & new_G1055_ & new_G1038_ & new_G1093_;
  assign new_G1125_ = new_G1026_ & new_G1050_;
  assign new_G1126_ = new_G1068_ & new_G1038_ & new_G1026_;
  assign new_G1127_ = new_G1038_ & new_G1086_ & new_G1055_ & new_G1026_;
  assign new_G1128_ = new_G1038_ & new_G1102_ & new_G1026_ & new_G1074_ & new_G1055_;
  assign new_G1132_ = new_G1038_ & new_G1068_;
  assign new_G1133_ = new_G1038_ & new_G1055_ & new_G1086_;
  assign new_G1134_ = new_G1038_ & new_G1102_ & new_G1074_ & new_G1055_;
  assign new_G1137_ = new_G1086_ & new_G1055_;
  assign new_G1138_ = new_G1102_ & new_G1074_ & new_G1055_;
  assign new_G1141_ = new_G1074_ & new_G1102_;
  assign new_G1221_ = ~new_G1217_;
  assign new_G1230_ = ~new_G1226_;
  assign new_G1244_ = ~new_G1240_;
  assign new_G1253_ = ~new_G1249_;
  assign new_G1267_ = ~new_G1263_;
  assign new_G1276_ = ~new_G1272_;
  assign new_G1284_ = new_G1235_;
  assign new_G1288_ = new_G1235_;
  assign new_G1292_ = new_G1258_;
  assign new_G1296_ = new_G1258_;
  assign new_G1300_ = new_G1281_;
  assign new_G1304_ = new_G1281_;
  assign new_G1702_ = new_G1546_ & new_G1556_ & new_G1687_ & new_G1573_;
  assign new_G1705_ = new_G1546_ & new_G1567_;
  assign new_G1706_ = new_G1584_ & new_G1556_ & new_G1546_;
  assign new_G1707_ = new_G1556_ & new_G1590_ & new_G1573_ & new_G1546_;
  assign new_G1709_ = new_G1556_ & new_G1584_;
  assign new_G1710_ = new_G1556_ & new_G1573_ & new_G1590_;
  assign new_G1711_ = new_G1556_ & new_G1687_ & new_G1573_;
  assign new_G1712_ = new_G1556_ & new_G1584_;
  assign new_G1713_ = new_G1556_ & new_G1573_ & new_G1590_;
  assign new_G1714_ = new_G1573_ & new_G1590_;
  assign new_G1718_ = new_G1598_ & new_G1609_ & new_G1630_ & new_G1695_ & new_G1655_;
  assign new_G1722_ = new_G1598_ & new_G1624_;
  assign new_G1723_ = new_G1647_ & new_G1609_ & new_G1598_;
  assign new_G1724_ = new_G1609_ & new_G1669_ & new_G1630_ & new_G1598_;
  assign new_G1725_ = new_G1609_ & new_G1677_ & new_G1598_ & new_G1655_ & new_G1630_;
  assign new_G1733_ = new_G1609_ & new_G1647_;
  assign new_G1734_ = new_G1609_ & new_G1630_ & new_G1669_;
  assign new_G1735_ = new_G1609_ & new_G1677_ & new_G1655_ & new_G1630_;
  assign new_G1736_ = new_G1655_ & new_G1609_ & new_G1695_ & new_G1630_;
  assign new_G1737_ = new_G1609_ & new_G1647_;
  assign new_G1738_ = new_G1609_ & new_G1630_ & new_G1669_;
  assign new_G1739_ = new_G1609_ & new_G1677_ & new_G1655_ & new_G1630_;
  assign new_G1740_ = new_G1630_ & new_G1669_;
  assign new_G1741_ = new_G1677_ & new_G1655_ & new_G1630_;
  assign new_G1742_ = new_G1655_ & new_G1695_ & new_G1630_;
  assign new_G1743_ = new_G1630_ & new_G1669_;
  assign new_G1744_ = new_G1677_ & new_G1655_ & new_G1630_;
  assign new_G1745_ = new_G1655_ & new_G1677_;
  assign new_G1749_ = new_G1687_ & new_G1573_;
  assign new_G1750_ = new_G1695_ & new_G1655_;
  assign new_G1935_ = new_G1795_ & new_G1822_ & new_G1805_ & new_G1850_;
  assign new_G1938_ = new_G1795_ & new_G1816_;
  assign new_G1939_ = new_G1834_ & new_G1805_ & new_G1795_;
  assign new_G1940_ = new_G1805_ & new_G1841_ & new_G1822_ & new_G1795_;
  assign new_G1942_ = new_G1805_ & new_G1834_;
  assign new_G1943_ = new_G1805_ & new_G1822_ & new_G1841_;
  assign new_G1944_ = new_G1805_ & new_G1850_ & new_G1822_;
  assign new_G1945_ = new_G1805_ & new_G1834_;
  assign new_G1946_ = new_G1805_ & new_G1841_ & new_G1822_;
  assign new_G1947_ = new_G1822_ & new_G1841_;
  assign new_G1948_ = new_G1850_ & new_G1822_;
  assign new_G1949_ = new_G1822_ & new_G1841_;
  assign new_G1950_ = new_G1903_ & new_G1859_ & new_G1885_ & new_G1869_ & new_G1921_;
  assign new_G1953_ = new_G1859_ & new_G1880_;
  assign new_G1954_ = new_G1897_ & new_G1869_ & new_G1859_;
  assign new_G1955_ = new_G1869_ & new_G1914_ & new_G1885_ & new_G1859_;
  assign new_G1956_ = new_G1869_ & new_G1929_ & new_G1859_ & new_G1903_ & new_G1885_;
  assign new_G1960_ = new_G1869_ & new_G1897_;
  assign new_G1961_ = new_G1869_ & new_G1885_ & new_G1914_;
  assign new_G1962_ = new_G1869_ & new_G1929_ & new_G1903_ & new_G1885_;
  assign new_G1965_ = new_G1914_ & new_G1885_;
  assign new_G1966_ = new_G1929_ & new_G1903_ & new_G1885_;
  assign new_G1969_ = new_G1903_ & new_G1929_;
  assign new_G2343_ = ~new_G2341_ | ~new_G2342_;
  assign new_G2354_ = ~new_G2352_ | ~new_G2353_;
  assign new_G2372_ = ~new_G2370_ | ~new_G2371_;
  assign new_G2400_ = ~new_G2398_ | ~new_G2399_;
  assign new_G2409_ = ~new_G2407_ | ~new_G2408_;
  assign new_G2420_ = ~new_G2418_ | ~new_G2419_;
  assign new_G2436_ = ~new_G2434_ | ~new_G2435_;
  assign new_G2454_ = ~new_G2452_ | ~new_G2453_;
  assign new_G2470_ = ~new_G5932_ | ~new_G5935_;
  assign new_G5936_ = ~new_G5932_;
  assign new_G5983_ = ~new_G5977_;
  assign new_G2589_ = ~new_G2587_ | ~new_G2588_;
  assign new_G2600_ = ~new_G2598_ | ~new_G2599_;
  assign new_G2618_ = ~new_G2616_ | ~new_G2617_;
  assign new_G2643_ = ~new_G2641_ | ~new_G2642_;
  assign new_G2655_ = ~new_G2653_ | ~new_G2654_;
  assign new_G2676_ = ~new_G2674_ | ~new_G2675_;
  assign new_G2701_ = ~new_G2699_ | ~new_G2700_;
  assign new_G2734_ = ~new_G2732_ | ~new_G2733_;
  assign new_G2740_ = ~new_G6052_ | ~new_G6055_;
  assign new_G6056_ = ~new_G6052_;
  assign new_G3022_ = new_G2956_ & new_G2965_ & new_G3018_ & new_G2973_;
  assign new_G3025_ = new_G2956_ & new_G2970_;
  assign new_G3026_ = new_G2977_ & new_G2965_ & new_G2956_;
  assign new_G3027_ = new_G2965_ & new_G2979_ & new_G2973_ & new_G2956_;
  assign new_G3029_ = new_G2982_ & new_G2992_ & new_G3001_ & new_G3021_ & new_G3009_;
  assign new_G3030_ = new_G2982_ & new_G2998_;
  assign new_G3031_ = new_G3006_ & new_G2992_ & new_G2982_;
  assign new_G3032_ = new_G2992_ & new_G3013_ & new_G3001_ & new_G2982_;
  assign new_G3033_ = new_G2992_ & new_G3015_ & new_G2982_ & new_G3009_ & new_G3001_;
  assign new_G3052_ = ~new_G3050_ | ~new_G3051_;
  assign new_G3062_ = ~new_G3060_ | ~new_G3061_;
  assign new_G3071_ = ~new_G3069_ | ~new_G3070_;
  assign new_G3082_ = ~new_G3080_ | ~new_G3081_;
  assign new_G3093_ = ~new_G3091_ | ~new_G3092_;
  assign new_G3102_ = ~new_G3100_ | ~new_G3101_;
  assign new_G3110_ = ~new_G3108_ | ~new_G3109_;
  assign new_G3119_ = ~new_G3117_ | ~new_G3118_;
  assign new_G3122_ = ~new_G3120_ | ~new_G3121_;
  assign new_G3228_ = new_G3176_ & new_G3186_ & new_G3195_ & new_G3215_ & new_G3203_;
  assign new_G3231_ = new_G3176_ & new_G3192_;
  assign new_G3232_ = new_G3200_ & new_G3186_ & new_G3176_;
  assign new_G3233_ = new_G3186_ & new_G3207_ & new_G3195_ & new_G3176_;
  assign new_G3234_ = new_G3186_ & new_G3209_ & new_G3176_ & new_G3203_ & new_G3195_;
  assign new_G3283_ = ~new_G3281_ | ~new_G3282_;
  assign new_G3295_ = ~new_G3293_ | ~new_G3294_;
  assign new_G3314_ = ~new_G3312_ | ~new_G3313_;
  assign new_G3344_ = ~new_G3342_ | ~new_G3343_;
  assign new_G3353_ = ~new_G3351_ | ~new_G3352_;
  assign new_G3365_ = ~new_G3363_ | ~new_G3364_;
  assign new_G3381_ = ~new_G3379_ | ~new_G3380_;
  assign new_G3399_ = ~new_G3397_ | ~new_G3398_;
  assign new_G3417_ = ~new_G3415_ | ~new_G3416_;
  assign new_G6685_ = ~new_G6679_;
  assign new_G3508_ = ~new_G3504_;
  assign new_G3517_ = ~new_G3513_;
  assign new_G3527_ = ~new_G3525_ | ~new_G3526_;
  assign new_G3536_ = ~new_G3534_ | ~new_G3535_;
  assign new_G3545_ = ~new_G3543_ | ~new_G3544_;
  assign new_G3550_ = ~new_G3548_ | ~new_G3549_;
  assign new_G3559_ = ~new_G3557_ | ~new_G3558_;
  assign new_G3568_ = ~new_G3566_ | ~new_G3567_;
  assign new_G3571_ = new_G3522_;
  assign new_G3575_ = new_G3522_;
  assign new_G3845_ = ~new_G3843_ | ~new_G3844_;
  assign new_G3856_ = ~new_G3854_ | ~new_G3855_;
  assign new_G3874_ = ~new_G3872_ | ~new_G3873_;
  assign new_G3899_ = ~new_G3897_ | ~new_G3898_;
  assign new_G3911_ = ~new_G3909_ | ~new_G3910_;
  assign new_G3932_ = ~new_G3930_ | ~new_G3931_;
  assign new_G3957_ = ~new_G3955_ | ~new_G3956_;
  assign new_G3989_ = ~new_G3987_ | ~new_G3988_;
  assign new_G3997_ = ~new_G3995_ | ~new_G3996_;
  assign new_G4180_ = ~new_G4178_ | ~new_G4179_;
  assign new_G4189_ = ~new_G4187_ | ~new_G4188_;
  assign new_G4198_ = ~new_G4196_ | ~new_G4197_;
  assign new_G4207_ = ~new_G4203_;
  assign new_G4216_ = ~new_G4212_;
  assign new_G4221_ = ~new_G4219_ | ~new_G4220_;
  assign new_G4230_ = ~new_G4226_;
  assign new_G4239_ = ~new_G4235_;
  assign new_G4263_ = new_G4244_;
  assign new_G4267_ = new_G4244_;
  assign new_G4291_ = ~new_G4289_ | ~new_G4290_;
  assign new_G4300_ = ~new_G4298_ | ~new_G4299_;
  assign new_G4308_ = ~new_G4306_ | ~new_G4307_;
  assign new_G4317_ = ~new_G4315_ | ~new_G4316_;
  assign new_G4327_ = ~new_G4325_ | ~new_G4326_;
  assign new_G4336_ = ~new_G4334_ | ~new_G4335_;
  assign new_G4344_ = ~new_G4342_ | ~new_G4343_;
  assign new_G4352_ = ~new_G4350_ | ~new_G4351_;
  assign new_G4355_ = ~new_G4353_ | ~new_G4354_;
  assign new_G4535_ = ~new_G4531_;
  assign new_G4544_ = ~new_G4540_;
  assign new_G4558_ = ~new_G4554_;
  assign new_G4563_ = ~new_G4561_ | ~new_G4562_;
  assign new_G4572_ = ~new_G4570_ | ~new_G4571_;
  assign new_G4577_ = ~new_G4575_ | ~new_G4576_;
  assign new_G4586_ = ~new_G4584_ | ~new_G4585_;
  assign new_G4595_ = ~new_G4593_ | ~new_G4594_;
  assign new_G4598_ = new_G4549_;
  assign new_G4602_ = new_G4549_;
  assign new_G4716_ = new_G1921_;
  assign new_G4724_ = new_G1859_;
  assign new_G4732_ = new_G1869_;
  assign new_G4740_ = new_G1885_;
  assign new_G4748_ = new_G1903_;
  assign new_G4756_ = new_G1093_;
  assign new_G4764_ = new_G1026_;
  assign new_G4772_ = new_G1038_;
  assign new_G4780_ = new_G1055_;
  assign new_G4788_ = new_G1074_;
  assign new_G4939_ = ~new_G4937_ | ~new_G4938_;
  assign new_G4980_ = ~new_G4978_ | ~new_G4979_;
  assign new_G5044_ = new_G895_;
  assign new_G5054_ = new_G853_;
  assign new_G5064_ = new_G792_;
  assign new_G5074_ = new_G827_;
  assign new_G5084_ = new_G805_;
  assign new_G5094_ = new_G805_;
  assign new_G5132_ = new_G895_;
  assign new_G5142_ = new_G853_;
  assign new_G5152_ = new_G792_;
  assign new_G5162_ = new_G827_;
  assign new_G5365_ = ~new_G5359_;
  assign new_G5366_ = ~new_G5362_;
  assign new_G5488_ = new_G1687_;
  assign new_G5498_ = new_G1573_;
  assign new_G5508_ = new_G1546_;
  assign new_G5518_ = new_G1556_;
  assign new_G5546_ = new_G1687_;
  assign new_G5556_ = new_G1573_;
  assign new_G5566_ = new_G1546_;
  assign new_G5576_ = new_G1556_;
  assign new_G5614_ = new_G1695_;
  assign new_G5624_ = new_G1655_;
  assign new_G5634_ = new_G1598_;
  assign new_G5644_ = new_G1630_;
  assign new_G5654_ = new_G1609_;
  assign new_G5664_ = new_G1609_;
  assign new_G5702_ = new_G1695_;
  assign new_G5712_ = new_G1655_;
  assign new_G5722_ = new_G1598_;
  assign new_G5732_ = new_G1630_;
  assign new_G5820_ = new_G1795_;
  assign new_G5828_ = new_G1795_;
  assign new_G5836_ = new_G1805_;
  assign new_G5844_ = new_G1805_;
  assign new_G5852_ = new_G1822_;
  assign new_G5860_ = new_G1822_;
  assign new_G6121_ = ~new_G6115_;
  assign new_G6179_ = ~new_G6173_;
  assign new_G6261_ = new_G2724_;
  assign new_G7359_ = ~new_G7353_;
  assign new_G7360_ = ~new_G7356_;
  assign new_G7343_ = ~new_G7337_;
  assign new_G7344_ = ~new_G7340_;
  assign new_G6809_ = ~new_G6763_ | ~new_G6764_;
  assign new_G6812_ = ~new_G6753_ | ~new_G6754_;
  assign new_G6819_ = ~new_G6807_ | ~new_G6808_;
  assign new_G6822_ = ~new_G6797_ | ~new_G6798_;
  assign new_G6989_ = ~new_G6983_;
  assign new_G7135_ = ~new_G7129_;
  assign new_G7345_ = ~new_G7291_ | ~new_G7292_;
  assign new_G7348_ = ~new_G7281_ | ~new_G7282_;
  assign new_G7601_ = ~new_G7595_;
  assign new_G7602_ = ~new_G7598_;
  assign new_G7603_ = ~new_G7549_ | ~new_G7550_;
  assign new_G7606_ = ~new_G7539_ | ~new_G7540_;
  assign new_G7611_ = ~new_G7593_ | ~new_G7594_;
  assign new_G7614_ = ~new_G7583_ | ~new_G7584_;
  assign new_G929_ = new_G928_ | new_G927_ | new_G926_ | new_G802_ | new_G925_;
  assign new_G950_ = new_G868_ | new_G949_;
  assign new_G1129_ = new_G1128_ | new_G1127_ | new_G1126_ | new_G1035_ | new_G1125_;
  assign new_G1708_ = new_G1707_ | new_G1706_ | new_G1553_ | new_G1705_;
  assign new_G1715_ = new_G1584_ | new_G1714_;
  assign new_G1726_ = new_G1725_ | new_G1724_ | new_G1723_ | new_G1606_ | new_G1722_;
  assign new_G1746_ = new_G1669_ | new_G1745_;
  assign new_G1941_ = new_G1940_ | new_G1939_ | new_G1802_ | new_G1938_;
  assign new_G1957_ = new_G1956_ | new_G1955_ | new_G1954_ | new_G1866_ | new_G1953_;
  assign new_G2471_ = ~new_G5929_ | ~new_G5936_;
  assign new_G2741_ = ~new_G6049_ | ~new_G6056_;
  assign new_G3028_ = new_G3027_ | new_G3026_ | new_G2962_ | new_G3025_;
  assign new_G3034_ = new_G3033_ | new_G3032_ | new_G3031_ | new_G2989_ | new_G3030_;
  assign new_G3235_ = new_G3234_ | new_G3233_ | new_G3232_ | new_G3183_ | new_G3231_;
  assign new_G5014_ = new_G946_ | new_G945_ | new_G845_ | new_G944_;
  assign new_G5034_ = new_G940_ | new_G939_ | new_G938_ | new_G821_ | new_G937_;
  assign new_G5102_ = ~new_G948_ & ~new_G845_ & ~new_G947_;
  assign new_G5122_ = ~new_G943_ & ~new_G942_ & ~new_G821_ & ~new_G941_;
  assign new_G5367_ = ~new_G5362_ | ~new_G5365_;
  assign new_G5368_ = ~new_G5359_ | ~new_G5366_;
  assign new_G5478_ = new_G1711_ | new_G1710_ | new_G1567_ | new_G1709_;
  assign new_G5536_ = ~new_G1713_ & ~new_G1567_ & ~new_G1712_;
  assign new_G5584_ = new_G1742_ | new_G1741_ | new_G1647_ | new_G1740_;
  assign new_G5604_ = new_G1736_ | new_G1735_ | new_G1734_ | new_G1624_ | new_G1733_;
  assign new_G5672_ = ~new_G1744_ & ~new_G1647_ & ~new_G1743_;
  assign new_G5692_ = ~new_G1739_ & ~new_G1738_ & ~new_G1624_ & ~new_G1737_;
  assign new_G5817_ = new_G1944_ | new_G1943_ | new_G1816_ | new_G1942_;
  assign new_G5825_ = ~new_G1946_ & ~new_G1816_ & ~new_G1945_;
  assign new_G5833_ = new_G1948_ | new_G1834_ | new_G1947_;
  assign new_G5841_ = ~new_G1834_ & ~new_G1949_;
  assign new_G6340_ = ~new_G7356_ | ~new_G7359_;
  assign new_G6341_ = ~new_G7353_ | ~new_G7360_;
  assign new_G6350_ = ~new_G7340_ | ~new_G7343_;
  assign new_G6351_ = ~new_G7337_ | ~new_G7344_;
  assign new_G7436_ = ~new_G7598_ | ~new_G7601_;
  assign new_G7437_ = ~new_G7595_ | ~new_G7602_;
  assign new_G4720_ = ~new_G4716_;
  assign new_G4728_ = ~new_G4724_;
  assign new_G4736_ = ~new_G4732_;
  assign new_G4744_ = ~new_G4740_;
  assign new_G4752_ = ~new_G4748_;
  assign new_G4760_ = ~new_G4756_;
  assign new_G4768_ = ~new_G4764_;
  assign new_G4776_ = ~new_G4772_;
  assign new_G4784_ = ~new_G4780_;
  assign new_G4792_ = ~new_G4788_;
  assign new_G3350_ = ~new_G3344_;
  assign new_G2406_ = ~new_G2400_;
  assign new_G924_ = ~new_G920_;
  assign new_G5088_ = ~new_G5084_;
  assign new_G5098_ = ~new_G5094_;
  assign new_G997_ = new_G902_ & new_G920_;
  assign new_G1146_ = new_G1108_ & new_G1122_;
  assign new_G1287_ = ~new_G1284_;
  assign new_G1291_ = ~new_G1288_;
  assign new_G1295_ = ~new_G1292_;
  assign new_G1299_ = ~new_G1296_;
  assign new_G1303_ = ~new_G1300_;
  assign new_G1307_ = ~new_G1304_;
  assign new_G1309_ = new_G1284_ & new_G1226_ & new_G1217_;
  assign new_G1312_ = new_G1288_ & new_G1230_ & new_G1221_;
  assign new_G1315_ = new_G1292_ & new_G1249_ & new_G1240_;
  assign new_G1318_ = new_G1296_ & new_G1253_ & new_G1244_;
  assign new_G1321_ = new_G1300_ & new_G1272_ & new_G1263_;
  assign new_G1324_ = new_G1304_ & new_G1276_ & new_G1267_;
  assign new_G1721_ = ~new_G1718_;
  assign new_G5522_ = ~new_G5518_;
  assign new_G5580_ = ~new_G5576_;
  assign new_G5658_ = ~new_G5654_;
  assign new_G5668_ = ~new_G5664_;
  assign new_G1788_ = new_G1702_ & new_G1718_;
  assign new_G1974_ = new_G1935_ & new_G1950_;
  assign new_G5824_ = ~new_G5820_;
  assign new_G5832_ = ~new_G5828_;
  assign new_G5840_ = ~new_G5836_;
  assign new_G5848_ = ~new_G5844_;
  assign new_G1999_ = ~new_G5852_ | ~new_G5855_;
  assign new_G5856_ = ~new_G5852_;
  assign new_G2003_ = ~new_G5860_ | ~new_G5863_;
  assign new_G5864_ = ~new_G5860_;
  assign new_G2472_ = ~new_G2470_ | ~new_G2471_;
  assign new_G2487_ = new_G2343_ & new_G2372_ & new_G2354_ & new_G2400_;
  assign new_G2492_ = new_G2343_ & new_G2366_;
  assign new_G2493_ = new_G2384_ & new_G2354_ & new_G2343_;
  assign new_G2494_ = new_G2354_ & new_G2391_ & new_G2372_ & new_G2343_;
  assign new_G2500_ = new_G2354_ & new_G2384_;
  assign new_G2501_ = new_G2354_ & new_G2372_ & new_G2391_;
  assign new_G2502_ = new_G2354_ & new_G2400_ & new_G2372_;
  assign new_G2503_ = new_G2354_ & new_G2384_;
  assign new_G2504_ = new_G2354_ & new_G2391_ & new_G2372_;
  assign new_G2505_ = new_G2372_ & new_G2391_;
  assign new_G2506_ = new_G2400_ & new_G2372_;
  assign new_G2507_ = new_G2372_ & new_G2391_;
  assign new_G2511_ = new_G2409_ & new_G2431_;
  assign new_G2512_ = new_G2448_ & new_G2420_ & new_G2409_;
  assign new_G2513_ = new_G2420_ & new_G2465_ & new_G2436_ & new_G2409_;
  assign new_G2514_ = new_G2420_ & new_G2481_ & new_G2409_ & new_G2454_ & new_G2436_;
  assign new_G2518_ = new_G2420_ & new_G2448_;
  assign new_G2519_ = new_G2420_ & new_G2436_ & new_G2465_;
  assign new_G2520_ = new_G2420_ & new_G2481_ & new_G2454_ & new_G2436_;
  assign new_G2523_ = new_G2465_ & new_G2436_;
  assign new_G2524_ = new_G2481_ & new_G2454_ & new_G2436_;
  assign new_G2527_ = new_G2454_ & new_G2481_;
  assign new_G2742_ = ~new_G2740_ | ~new_G2741_;
  assign new_G2749_ = new_G2589_ & new_G2600_ & new_G2734_ & new_G2618_;
  assign new_G2754_ = new_G2589_ & new_G2612_;
  assign new_G2755_ = new_G2629_ & new_G2600_ & new_G2589_;
  assign new_G2756_ = new_G2600_ & new_G2635_ & new_G2618_ & new_G2589_;
  assign new_G2762_ = new_G2600_ & new_G2629_;
  assign new_G2763_ = new_G2600_ & new_G2618_ & new_G2635_;
  assign new_G2764_ = new_G2600_ & new_G2734_ & new_G2618_;
  assign new_G2765_ = new_G2600_ & new_G2629_;
  assign new_G2766_ = new_G2600_ & new_G2618_ & new_G2635_;
  assign new_G2767_ = new_G2618_ & new_G2635_;
  assign new_G2776_ = new_G2643_ & new_G2670_;
  assign new_G2777_ = new_G2693_ & new_G2655_ & new_G2643_;
  assign new_G2778_ = new_G2655_ & new_G2715_ & new_G2676_ & new_G2643_;
  assign new_G2779_ = new_G2655_ & new_G2724_ & new_G2643_ & new_G2701_ & new_G2676_;
  assign new_G2788_ = new_G2655_ & new_G2693_;
  assign new_G2789_ = new_G2655_ & new_G2676_ & new_G2715_;
  assign new_G2790_ = new_G2655_ & new_G2724_ & new_G2701_ & new_G2676_;
  assign new_G2792_ = new_G2655_ & new_G2693_;
  assign new_G2793_ = new_G2655_ & new_G2676_ & new_G2715_;
  assign new_G2794_ = new_G2655_ & new_G2724_ & new_G2701_ & new_G2676_;
  assign new_G2795_ = new_G2676_ & new_G2715_;
  assign new_G2796_ = new_G2724_ & new_G2701_ & new_G2676_;
  assign new_G2798_ = new_G2676_ & new_G2715_;
  assign new_G2799_ = new_G2724_ & new_G2701_ & new_G2676_;
  assign new_G2800_ = new_G2701_ & new_G2724_;
  assign new_G2804_ = new_G2734_ & new_G2618_;
  assign new_G3035_ = new_G3022_ & new_G3029_;
  assign new_G3045_ = new_G3022_ & new_G3034_;
  assign new_G3123_ = new_G3052_ & new_G3062_ & new_G3119_ & new_G3071_;
  assign new_G3128_ = new_G3052_ & new_G3068_;
  assign new_G3129_ = new_G3076_ & new_G3062_ & new_G3052_;
  assign new_G3130_ = new_G3062_ & new_G3079_ & new_G3071_ & new_G3052_;
  assign new_G3136_ = new_G3082_ & new_G3093_ & new_G3102_ & new_G3122_ & new_G3110_;
  assign new_G3139_ = new_G3082_ & new_G3099_;
  assign new_G3140_ = new_G3107_ & new_G3093_ & new_G3082_;
  assign new_G3141_ = new_G3093_ & new_G3114_ & new_G3102_ & new_G3082_;
  assign new_G3142_ = new_G3093_ & new_G3116_ & new_G3082_ & new_G3110_ & new_G3102_;
  assign new_G3249_ = new_G3216_ & new_G3228_;
  assign new_G3431_ = new_G3283_ & new_G3314_ & new_G3295_ & new_G3344_;
  assign new_G3434_ = new_G3283_ & new_G3308_;
  assign new_G3435_ = new_G3327_ & new_G3295_ & new_G3283_;
  assign new_G3436_ = new_G3295_ & new_G3335_ & new_G3314_ & new_G3283_;
  assign new_G3438_ = new_G3295_ & new_G3327_;
  assign new_G3439_ = new_G3295_ & new_G3314_ & new_G3335_;
  assign new_G3440_ = new_G3295_ & new_G3344_ & new_G3314_;
  assign new_G3441_ = new_G3295_ & new_G3327_;
  assign new_G3442_ = new_G3295_ & new_G3335_ & new_G3314_;
  assign new_G3443_ = new_G3314_ & new_G3335_;
  assign new_G3444_ = new_G3344_ & new_G3314_;
  assign new_G3445_ = new_G3314_ & new_G3335_;
  assign new_G3446_ = new_G3399_ & new_G3353_ & new_G3381_ & new_G3365_ & new_G3417_;
  assign new_G3449_ = new_G3353_ & new_G3376_;
  assign new_G3450_ = new_G3393_ & new_G3365_ & new_G3353_;
  assign new_G3451_ = new_G3365_ & new_G3410_ & new_G3381_ & new_G3353_;
  assign new_G3452_ = new_G3365_ & new_G3425_ & new_G3353_ & new_G3399_ & new_G3381_;
  assign new_G3456_ = new_G3365_ & new_G3393_;
  assign new_G3457_ = new_G3365_ & new_G3381_ & new_G3410_;
  assign new_G3458_ = new_G3365_ & new_G3425_ & new_G3399_ & new_G3381_;
  assign new_G3460_ = new_G3410_ & new_G3381_;
  assign new_G3461_ = new_G3425_ & new_G3399_ & new_G3381_;
  assign new_G3463_ = new_G3399_ & new_G3425_;
  assign new_G3531_ = ~new_G3527_;
  assign new_G3540_ = ~new_G3536_;
  assign new_G3554_ = ~new_G3550_;
  assign new_G3563_ = ~new_G3559_;
  assign new_G3574_ = ~new_G3571_;
  assign new_G3578_ = ~new_G3575_;
  assign new_G3579_ = new_G3545_;
  assign new_G3583_ = new_G3545_;
  assign new_G3587_ = new_G3568_;
  assign new_G3591_ = new_G3568_;
  assign new_G3596_ = new_G3571_ & new_G3513_ & new_G3504_;
  assign new_G3599_ = new_G3575_ & new_G3517_ & new_G3508_;
  assign new_G4004_ = new_G3845_ & new_G3856_ & new_G3989_ & new_G3874_;
  assign new_G4007_ = new_G3845_ & new_G3868_;
  assign new_G4008_ = new_G3885_ & new_G3856_ & new_G3845_;
  assign new_G4009_ = new_G3856_ & new_G3891_ & new_G3874_ & new_G3845_;
  assign new_G4011_ = new_G3856_ & new_G3885_;
  assign new_G4012_ = new_G3856_ & new_G3874_ & new_G3891_;
  assign new_G4013_ = new_G3856_ & new_G3989_ & new_G3874_;
  assign new_G4014_ = new_G3856_ & new_G3885_;
  assign new_G4015_ = new_G3856_ & new_G3874_ & new_G3891_;
  assign new_G4016_ = new_G3874_ & new_G3891_;
  assign new_G4020_ = new_G3899_ & new_G3911_ & new_G3932_ & new_G3997_ & new_G3957_;
  assign new_G4024_ = new_G3899_ & new_G3926_;
  assign new_G4025_ = new_G3949_ & new_G3911_ & new_G3899_;
  assign new_G4026_ = new_G3911_ & new_G3971_ & new_G3932_ & new_G3899_;
  assign new_G4027_ = new_G3911_ & new_G3979_ & new_G3899_ & new_G3957_ & new_G3932_;
  assign new_G4035_ = new_G3911_ & new_G3949_;
  assign new_G4036_ = new_G3911_ & new_G3932_ & new_G3971_;
  assign new_G4037_ = new_G3911_ & new_G3979_ & new_G3957_ & new_G3932_;
  assign new_G4038_ = new_G3957_ & new_G3911_ & new_G3997_ & new_G3932_;
  assign new_G4039_ = new_G3911_ & new_G3949_;
  assign new_G4040_ = new_G3911_ & new_G3932_ & new_G3971_;
  assign new_G4041_ = new_G3911_ & new_G3979_ & new_G3957_ & new_G3932_;
  assign new_G4042_ = new_G3932_ & new_G3971_;
  assign new_G4043_ = new_G3979_ & new_G3957_ & new_G3932_;
  assign new_G4044_ = new_G3957_ & new_G3997_ & new_G3932_;
  assign new_G4045_ = new_G3932_ & new_G3971_;
  assign new_G4046_ = new_G3979_ & new_G3957_ & new_G3932_;
  assign new_G4047_ = new_G3957_ & new_G3979_;
  assign new_G4051_ = new_G3989_ & new_G3874_;
  assign new_G4052_ = new_G3997_ & new_G3957_;
  assign new_G4184_ = ~new_G4180_;
  assign new_G4193_ = ~new_G4189_;
  assign new_G4247_ = new_G4198_;
  assign new_G4251_ = new_G4198_;
  assign new_G4255_ = new_G4221_;
  assign new_G4259_ = new_G4221_;
  assign new_G4266_ = ~new_G4263_;
  assign new_G4270_ = ~new_G4267_;
  assign new_G4284_ = new_G4263_ & new_G4235_ & new_G4226_;
  assign new_G4287_ = new_G4267_ & new_G4239_ & new_G4230_;
  assign new_G4356_ = new_G4291_ & new_G4300_ & new_G4352_ & new_G4308_;
  assign new_G4361_ = new_G4291_ & new_G4305_;
  assign new_G4362_ = new_G4312_ & new_G4300_ & new_G4291_;
  assign new_G4363_ = new_G4300_ & new_G4314_ & new_G4308_ & new_G4291_;
  assign new_G4369_ = new_G4317_ & new_G4327_ & new_G4336_ & new_G4355_ & new_G4344_;
  assign new_G4372_ = new_G4317_ & new_G4333_;
  assign new_G4373_ = new_G4341_ & new_G4327_ & new_G4317_;
  assign new_G4374_ = new_G4327_ & new_G4348_ & new_G4336_ & new_G4317_;
  assign new_G4375_ = new_G4327_ & new_G4349_ & new_G4317_ & new_G4344_ & new_G4336_;
  assign new_G4567_ = ~new_G4563_;
  assign new_G4581_ = ~new_G4577_;
  assign new_G4590_ = ~new_G4586_;
  assign new_G4601_ = ~new_G4598_;
  assign new_G4605_ = ~new_G4602_;
  assign new_G4606_ = new_G4572_;
  assign new_G4610_ = new_G4572_;
  assign new_G4614_ = new_G4595_;
  assign new_G4618_ = new_G4595_;
  assign new_G4623_ = new_G4598_ & new_G4540_ & new_G4531_;
  assign new_G4626_ = new_G4602_ & new_G4544_ & new_G4535_;
  assign new_G4796_ = new_G3417_;
  assign new_G4804_ = new_G3353_;
  assign new_G4812_ = new_G3365_;
  assign new_G4820_ = new_G3381_;
  assign new_G4828_ = new_G3399_;
  assign new_G4844_ = new_G2409_;
  assign new_G4852_ = new_G2420_;
  assign new_G4860_ = new_G2436_;
  assign new_G4868_ = new_G2454_;
  assign new_G4945_ = ~new_G4939_;
  assign new_G4948_ = ~new_G4939_ | ~new_G4946_;
  assign new_G4986_ = ~new_G4980_;
  assign new_G4989_ = ~new_G4980_ | ~new_G4987_;
  assign new_G5048_ = ~new_G5044_;
  assign new_G5058_ = ~new_G5054_;
  assign new_G5068_ = ~new_G5064_;
  assign new_G5078_ = ~new_G5074_;
  assign new_G5166_ = ~new_G5162_;
  assign new_G5136_ = ~new_G5132_;
  assign new_G5146_ = ~new_G5142_;
  assign new_G5156_ = ~new_G5152_;
  assign new_G5388_ = ~new_G5367_ | ~new_G5368_;
  assign new_G5492_ = ~new_G5488_;
  assign new_G5502_ = ~new_G5498_;
  assign new_G5512_ = ~new_G5508_;
  assign new_G5550_ = ~new_G5546_;
  assign new_G5560_ = ~new_G5556_;
  assign new_G5570_ = ~new_G5566_;
  assign new_G5618_ = ~new_G5614_;
  assign new_G5628_ = ~new_G5624_;
  assign new_G5638_ = ~new_G5634_;
  assign new_G5648_ = ~new_G5644_;
  assign new_G5736_ = ~new_G5732_;
  assign new_G5706_ = ~new_G5702_;
  assign new_G5716_ = ~new_G5712_;
  assign new_G5726_ = ~new_G5722_;
  assign new_G5940_ = new_G2343_;
  assign new_G5948_ = new_G2343_;
  assign new_G5956_ = new_G2354_;
  assign new_G5964_ = new_G2354_;
  assign new_G5972_ = new_G2372_;
  assign new_G5980_ = new_G2372_;
  assign new_G6080_ = new_G2734_;
  assign new_G6090_ = new_G2618_;
  assign new_G6100_ = new_G2589_;
  assign new_G6110_ = new_G2600_;
  assign new_G6138_ = new_G2734_;
  assign new_G6148_ = new_G2618_;
  assign new_G6158_ = new_G2589_;
  assign new_G6168_ = new_G2600_;
  assign new_G6216_ = new_G2701_;
  assign new_G6226_ = new_G2643_;
  assign new_G6236_ = new_G2676_;
  assign new_G6246_ = new_G2655_;
  assign new_G6256_ = new_G2655_;
  assign new_G6267_ = ~new_G6261_;
  assign new_G6304_ = new_G2701_;
  assign new_G6314_ = new_G2643_;
  assign new_G6324_ = new_G2676_;
  assign new_G6342_ = ~new_G6340_ | ~new_G6341_;
  assign new_G6352_ = ~new_G6350_ | ~new_G6351_;
  assign new_G7351_ = ~new_G7345_;
  assign new_G7352_ = ~new_G7348_;
  assign new_G6642_ = new_G3283_;
  assign new_G6650_ = new_G3283_;
  assign new_G6658_ = new_G3295_;
  assign new_G6666_ = new_G3295_;
  assign new_G6674_ = new_G3314_;
  assign new_G6682_ = new_G3314_;
  assign new_G6815_ = ~new_G6809_;
  assign new_G6816_ = ~new_G6812_;
  assign new_G6825_ = ~new_G6819_;
  assign new_G6826_ = ~new_G6822_;
  assign new_G6948_ = new_G3989_;
  assign new_G6958_ = new_G3874_;
  assign new_G6968_ = new_G3845_;
  assign new_G6978_ = new_G3856_;
  assign new_G7006_ = new_G3989_;
  assign new_G7016_ = new_G3874_;
  assign new_G7026_ = new_G3845_;
  assign new_G7036_ = new_G3856_;
  assign new_G7074_ = new_G3997_;
  assign new_G7084_ = new_G3957_;
  assign new_G7094_ = new_G3899_;
  assign new_G7104_ = new_G3932_;
  assign new_G7114_ = new_G3911_;
  assign new_G7124_ = new_G3911_;
  assign new_G7162_ = new_G3997_;
  assign new_G7172_ = new_G3957_;
  assign new_G7182_ = new_G3899_;
  assign new_G7192_ = new_G3932_;
  assign new_G7438_ = ~new_G7436_ | ~new_G7437_;
  assign new_G7617_ = ~new_G7611_;
  assign new_G7618_ = ~new_G7614_;
  assign new_G7609_ = ~new_G7603_;
  assign new_G7610_ = ~new_G7606_;
  assign new_G1151_ = new_G1129_ & new_G1108_;
  assign new_G1002_ = new_G902_ & new_G929_;
  assign new_G933_ = ~new_G929_;
  assign new_G1308_ = new_G1287_ & new_G1221_ & new_G1226_;
  assign new_G1311_ = new_G1291_ & new_G1217_ & new_G1230_;
  assign new_G1314_ = new_G1295_ & new_G1244_ & new_G1249_;
  assign new_G1317_ = new_G1299_ & new_G1240_ & new_G1253_;
  assign new_G1320_ = new_G1303_ & new_G1267_ & new_G1272_;
  assign new_G1323_ = new_G1307_ & new_G1263_ & new_G1276_;
  assign new_G1730_ = ~new_G1726_;
  assign new_G1789_ = new_G1702_ & new_G1726_;
  assign new_G1981_ = new_G1957_ & new_G1935_;
  assign new_G5823_ = ~new_G5817_;
  assign new_G1986_ = ~new_G5817_ | ~new_G5824_;
  assign new_G5831_ = ~new_G5825_;
  assign new_G1989_ = ~new_G5825_ | ~new_G5832_;
  assign new_G5839_ = ~new_G5833_;
  assign new_G1993_ = ~new_G5833_ | ~new_G5840_;
  assign new_G5847_ = ~new_G5841_;
  assign new_G1996_ = ~new_G5841_ | ~new_G5848_;
  assign new_G2000_ = ~new_G5849_ | ~new_G5856_;
  assign new_G2004_ = ~new_G5857_ | ~new_G5864_;
  assign new_G2495_ = new_G2494_ | new_G2493_ | new_G2351_ | new_G2492_;
  assign new_G2515_ = new_G2514_ | new_G2513_ | new_G2512_ | new_G2417_ | new_G2511_;
  assign new_G2757_ = new_G2756_ | new_G2755_ | new_G2597_ | new_G2754_;
  assign new_G2768_ = new_G2629_ | new_G2767_;
  assign new_G2780_ = new_G2779_ | new_G2778_ | new_G2777_ | new_G2652_ | new_G2776_;
  assign new_G2801_ = new_G2715_ | new_G2800_;
  assign new_G3046_ = new_G3028_ | new_G3045_;
  assign new_G3131_ = new_G3130_ | new_G3129_ | new_G3059_ | new_G3128_;
  assign new_G3143_ = new_G3142_ | new_G3141_ | new_G3140_ | new_G3090_ | new_G3139_;
  assign new_G3238_ = ~new_G3235_;
  assign new_G3258_ = new_G3216_ & new_G3235_;
  assign new_G3437_ = new_G3436_ | new_G3435_ | new_G3292_ | new_G3434_;
  assign new_G3453_ = new_G3452_ | new_G3451_ | new_G3450_ | new_G3362_ | new_G3449_;
  assign new_G3595_ = new_G3574_ & new_G3508_ & new_G3513_;
  assign new_G3598_ = new_G3578_ & new_G3504_ & new_G3517_;
  assign new_G4010_ = new_G4009_ | new_G4008_ | new_G3853_ | new_G4007_;
  assign new_G4017_ = new_G3885_ | new_G4016_;
  assign new_G4028_ = new_G4027_ | new_G4026_ | new_G4025_ | new_G3908_ | new_G4024_;
  assign new_G4048_ = new_G3971_ | new_G4047_;
  assign new_G4283_ = new_G4266_ & new_G4230_ & new_G4235_;
  assign new_G4286_ = new_G4270_ & new_G4226_ & new_G4239_;
  assign new_G4364_ = new_G4363_ | new_G4362_ | new_G4297_ | new_G4361_;
  assign new_G4376_ = new_G4375_ | new_G4374_ | new_G4373_ | new_G4324_ | new_G4372_;
  assign new_G4622_ = new_G4601_ & new_G4535_ & new_G4540_;
  assign new_G4625_ = new_G4605_ & new_G4531_ & new_G4544_;
  assign new_G4947_ = ~new_G4942_ | ~new_G4945_;
  assign new_G4988_ = ~new_G4983_ | ~new_G4986_;
  assign new_G5018_ = ~new_G5014_;
  assign new_G5019_ = ~new_G5014_ | ~new_G5017_;
  assign new_G5024_ = new_G950_ | new_G956_;
  assign new_G5038_ = ~new_G5034_;
  assign new_G5106_ = ~new_G5102_;
  assign new_G5107_ = ~new_G5102_ | ~new_G5105_;
  assign new_G5112_ = ~new_G950_;
  assign new_G5126_ = ~new_G5122_;
  assign new_G5468_ = new_G1715_ | new_G1749_;
  assign new_G5482_ = ~new_G5478_;
  assign new_G5526_ = ~new_G1715_;
  assign new_G5540_ = ~new_G5536_;
  assign new_G5588_ = ~new_G5584_;
  assign new_G5589_ = ~new_G5584_ | ~new_G5587_;
  assign new_G5594_ = new_G1746_ | new_G1750_;
  assign new_G5608_ = ~new_G5604_;
  assign new_G5676_ = ~new_G5672_;
  assign new_G5677_ = ~new_G5672_ | ~new_G5675_;
  assign new_G5682_ = ~new_G1746_;
  assign new_G5696_ = ~new_G5692_;
  assign new_G5937_ = new_G2502_ | new_G2501_ | new_G2366_ | new_G2500_;
  assign new_G5945_ = ~new_G2504_ & ~new_G2366_ & ~new_G2503_;
  assign new_G5953_ = new_G2506_ | new_G2384_ | new_G2505_;
  assign new_G5961_ = ~new_G2384_ & ~new_G2507_;
  assign new_G6070_ = new_G2764_ | new_G2763_ | new_G2612_ | new_G2762_;
  assign new_G6128_ = ~new_G2766_ & ~new_G2612_ & ~new_G2765_;
  assign new_G6264_ = ~new_G2799_ & ~new_G2693_ & ~new_G2798_;
  assign new_G6284_ = ~new_G2794_ & ~new_G2793_ & ~new_G2670_ & ~new_G2792_;
  assign new_G6360_ = ~new_G7348_ | ~new_G7351_;
  assign new_G6361_ = ~new_G7345_ | ~new_G7352_;
  assign new_G6639_ = new_G3440_ | new_G3439_ | new_G3308_ | new_G3438_;
  assign new_G6647_ = ~new_G3442_ & ~new_G3308_ & ~new_G3441_;
  assign new_G6655_ = new_G3444_ | new_G3327_ | new_G3443_;
  assign new_G6663_ = ~new_G3327_ & ~new_G3445_;
  assign new_G6817_ = ~new_G6812_ | ~new_G6815_;
  assign new_G6818_ = ~new_G6809_ | ~new_G6816_;
  assign new_G6827_ = ~new_G6822_ | ~new_G6825_;
  assign new_G6828_ = ~new_G6819_ | ~new_G6826_;
  assign new_G6938_ = new_G4013_ | new_G4012_ | new_G3868_ | new_G4011_;
  assign new_G6996_ = ~new_G4015_ & ~new_G3868_ & ~new_G4014_;
  assign new_G7044_ = new_G4044_ | new_G4043_ | new_G3949_ | new_G4042_;
  assign new_G7064_ = new_G4038_ | new_G4037_ | new_G4036_ | new_G3926_ | new_G4035_;
  assign new_G7132_ = ~new_G4046_ & ~new_G3949_ & ~new_G4045_;
  assign new_G7152_ = ~new_G4041_ & ~new_G4040_ & ~new_G3926_ & ~new_G4039_;
  assign new_G7446_ = ~new_G7614_ | ~new_G7617_;
  assign new_G7447_ = ~new_G7611_ | ~new_G7618_;
  assign new_G7456_ = ~new_G7606_ | ~new_G7609_;
  assign new_G7457_ = ~new_G7603_ | ~new_G7610_;
  assign new_G241_ = new_G1117_ | new_G1151_;
  assign new_G265_ = new_G908_ | new_G1002_;
  assign new_G2005_ = ~new_G2003_ | ~new_G2004_;
  assign new_G4800_ = ~new_G4796_;
  assign new_G4808_ = ~new_G4804_;
  assign new_G4816_ = ~new_G4812_;
  assign new_G4824_ = ~new_G4820_;
  assign new_G4832_ = ~new_G4828_;
  assign new_G4848_ = ~new_G4844_;
  assign new_G4856_ = ~new_G4852_;
  assign new_G4864_ = ~new_G4860_;
  assign new_G4872_ = ~new_G4868_;
  assign new_G1310_ = ~new_G1308_ & ~new_G1309_;
  assign new_G1313_ = ~new_G1311_ & ~new_G1312_;
  assign new_G1316_ = ~new_G1314_ & ~new_G1315_;
  assign new_G1319_ = ~new_G1317_ & ~new_G1318_;
  assign new_G1322_ = ~new_G1320_ & ~new_G1321_;
  assign new_G1325_ = ~new_G1323_ & ~new_G1324_;
  assign new_G5392_ = ~new_G5388_;
  assign new_G1790_ = new_G1708_ | new_G1789_;
  assign new_G1982_ = new_G1941_ | new_G1981_;
  assign new_G1985_ = ~new_G5820_ | ~new_G5823_;
  assign new_G1988_ = ~new_G5828_ | ~new_G5831_;
  assign new_G1992_ = ~new_G5836_ | ~new_G5839_;
  assign new_G1995_ = ~new_G5844_ | ~new_G5847_;
  assign new_G2001_ = ~new_G1999_ | ~new_G2000_;
  assign new_G2491_ = ~new_G2487_;
  assign new_G2508_ = new_G2454_ & new_G2409_ & new_G2436_ & new_G2420_ & new_G2472_;
  assign new_G2522_ = new_G2420_ & new_G2454_ & new_G2436_ & G4526 & new_G2472_;
  assign new_G2526_ = new_G2454_ & new_G2436_ & G4526 & new_G2472_;
  assign new_G2529_ = new_G2454_ & G4526 & new_G2472_;
  assign new_G2531_ = G4526 & new_G2472_;
  assign new_G5944_ = ~new_G5940_;
  assign new_G5952_ = ~new_G5948_;
  assign new_G5960_ = ~new_G5956_;
  assign new_G5968_ = ~new_G5964_;
  assign new_G2555_ = ~new_G5972_ | ~new_G5975_;
  assign new_G5976_ = ~new_G5972_;
  assign new_G2559_ = ~new_G5980_ | ~new_G5983_;
  assign new_G5984_ = ~new_G5980_;
  assign new_G2753_ = ~new_G2749_;
  assign new_G2771_ = new_G2643_ & new_G2655_ & new_G2676_ & new_G2742_ & new_G2701_;
  assign new_G2791_ = new_G2701_ & new_G2655_ & new_G2742_ & new_G2676_;
  assign new_G2797_ = new_G2701_ & new_G2742_ & new_G2676_;
  assign new_G2807_ = new_G2742_ & new_G2701_;
  assign new_G6114_ = ~new_G6110_;
  assign new_G6172_ = ~new_G6168_;
  assign new_G6250_ = ~new_G6246_;
  assign new_G6260_ = ~new_G6256_;
  assign new_G6346_ = ~new_G6342_;
  assign new_G6356_ = ~new_G6352_;
  assign new_G3127_ = ~new_G3123_;
  assign new_G3156_ = new_G3123_ & new_G3136_;
  assign new_G3259_ = new_G3223_ | new_G3258_;
  assign new_G3466_ = new_G3431_ & new_G3446_;
  assign new_G6646_ = ~new_G6642_;
  assign new_G6654_ = ~new_G6650_;
  assign new_G6662_ = ~new_G6658_;
  assign new_G6670_ = ~new_G6666_;
  assign new_G3483_ = ~new_G6674_ | ~new_G6677_;
  assign new_G6678_ = ~new_G6674_;
  assign new_G3487_ = ~new_G6682_ | ~new_G6685_;
  assign new_G6686_ = ~new_G6682_;
  assign new_G3582_ = ~new_G3579_;
  assign new_G3586_ = ~new_G3583_;
  assign new_G3590_ = ~new_G3587_;
  assign new_G3594_ = ~new_G3591_;
  assign new_G3597_ = ~new_G3595_ & ~new_G3596_;
  assign new_G3600_ = ~new_G3598_ & ~new_G3599_;
  assign new_G3602_ = new_G3579_ & new_G3536_ & new_G3527_;
  assign new_G3605_ = new_G3583_ & new_G3540_ & new_G3531_;
  assign new_G3608_ = new_G3587_ & new_G3559_ & new_G3550_;
  assign new_G3611_ = new_G3591_ & new_G3563_ & new_G3554_;
  assign new_G4023_ = ~new_G4020_;
  assign new_G6982_ = ~new_G6978_;
  assign new_G7040_ = ~new_G7036_;
  assign new_G7118_ = ~new_G7114_;
  assign new_G7128_ = ~new_G7124_;
  assign new_G4089_ = new_G4004_ & new_G4020_;
  assign new_G4250_ = ~new_G4247_;
  assign new_G4254_ = ~new_G4251_;
  assign new_G4258_ = ~new_G4255_;
  assign new_G4262_ = ~new_G4259_;
  assign new_G4272_ = new_G4247_ & new_G4189_ & new_G4180_;
  assign new_G4275_ = new_G4251_ & new_G4193_ & new_G4184_;
  assign new_G4278_ = new_G4255_ & new_G4212_ & new_G4203_;
  assign new_G4281_ = new_G4259_ & new_G4216_ & new_G4207_;
  assign new_G4285_ = ~new_G4283_ & ~new_G4284_;
  assign new_G4288_ = ~new_G4286_ & ~new_G4287_;
  assign new_G4360_ = ~new_G4356_;
  assign new_G4380_ = ~new_G4369_ | ~G89;
  assign new_G4386_ = new_G4356_ & new_G4369_;
  assign new_G7442_ = ~new_G7438_;
  assign new_G4609_ = ~new_G4606_;
  assign new_G4613_ = ~new_G4610_;
  assign new_G4617_ = ~new_G4614_;
  assign new_G4621_ = ~new_G4618_;
  assign new_G4624_ = ~new_G4622_ & ~new_G4623_;
  assign new_G4627_ = ~new_G4625_ & ~new_G4626_;
  assign new_G4629_ = new_G4606_ & new_G4563_ & new_G4554_;
  assign new_G4632_ = new_G4610_ & new_G4567_ & new_G4558_;
  assign new_G4635_ = new_G4614_ & new_G4586_ & new_G4577_;
  assign new_G4638_ = new_G4618_ & new_G4590_ & new_G4581_;
  assign new_G4836_ = new_G2472_;
  assign new_G4949_ = ~new_G4947_ | ~new_G4948_;
  assign new_G4990_ = ~new_G4988_ | ~new_G4989_;
  assign new_G5020_ = ~new_G5011_ | ~new_G5018_;
  assign new_G5108_ = ~new_G5099_ | ~new_G5106_;
  assign new_G5590_ = ~new_G5581_ | ~new_G5588_;
  assign new_G5678_ = ~new_G5669_ | ~new_G5676_;
  assign new_G6084_ = ~new_G6080_;
  assign new_G6094_ = ~new_G6090_;
  assign new_G6104_ = ~new_G6100_;
  assign new_G6142_ = ~new_G6138_;
  assign new_G6152_ = ~new_G6148_;
  assign new_G6162_ = ~new_G6158_;
  assign new_G6206_ = new_G2742_;
  assign new_G6220_ = ~new_G6216_;
  assign new_G6230_ = ~new_G6226_;
  assign new_G6240_ = ~new_G6236_;
  assign new_G6328_ = ~new_G6324_;
  assign new_G6294_ = new_G2742_;
  assign new_G6308_ = ~new_G6304_;
  assign new_G6318_ = ~new_G6314_;
  assign new_G6362_ = ~new_G6360_ | ~new_G6361_;
  assign new_G6840_ = ~new_G6817_ | ~new_G6818_;
  assign new_G6848_ = ~new_G6827_ | ~new_G6828_;
  assign new_G6952_ = ~new_G6948_;
  assign new_G6962_ = ~new_G6958_;
  assign new_G6972_ = ~new_G6968_;
  assign new_G7010_ = ~new_G7006_;
  assign new_G7020_ = ~new_G7016_;
  assign new_G7030_ = ~new_G7026_;
  assign new_G7078_ = ~new_G7074_;
  assign new_G7088_ = ~new_G7084_;
  assign new_G7098_ = ~new_G7094_;
  assign new_G7108_ = ~new_G7104_;
  assign new_G7196_ = ~new_G7192_;
  assign new_G7166_ = ~new_G7162_;
  assign new_G7176_ = ~new_G7172_;
  assign new_G7186_ = ~new_G7182_;
  assign new_G7448_ = ~new_G7446_ | ~new_G7447_;
  assign new_G7458_ = ~new_G7456_ | ~new_G7457_;
  assign new_G254_ = new_G3046_ & new_G3249_;
  assign new_G260_ = new_G3046_ & new_G3249_;
  assign new_G1987_ = ~new_G1985_ | ~new_G1986_;
  assign new_G1994_ = ~new_G1992_ | ~new_G1993_;
  assign new_G2002_ = ~new_G2001_;
  assign new_G962_ = new_G933_ & new_G924_;
  assign new_G1751_ = new_G1730_ & new_G1721_;
  assign new_G1990_ = ~new_G1988_ | ~new_G1989_;
  assign new_G1997_ = ~new_G1995_ | ~new_G1996_;
  assign new_G2499_ = ~new_G2495_;
  assign new_G2536_ = new_G2515_ & new_G2487_;
  assign new_G5943_ = ~new_G5937_;
  assign new_G2542_ = ~new_G5937_ | ~new_G5944_;
  assign new_G5951_ = ~new_G5945_;
  assign new_G2545_ = ~new_G5945_ | ~new_G5952_;
  assign new_G5959_ = ~new_G5953_;
  assign new_G2549_ = ~new_G5953_ | ~new_G5960_;
  assign new_G5967_ = ~new_G5961_;
  assign new_G2552_ = ~new_G5961_ | ~new_G5968_;
  assign new_G2556_ = ~new_G5969_ | ~new_G5976_;
  assign new_G2560_ = ~new_G5977_ | ~new_G5984_;
  assign new_G2761_ = ~new_G2757_;
  assign new_G2784_ = ~new_G2780_;
  assign new_G2853_ = new_G2749_ & new_G2780_;
  assign new_G3135_ = ~new_G3131_;
  assign new_G3146_ = ~new_G3143_;
  assign new_G3163_ = new_G3123_ & new_G3143_;
  assign new_G3467_ = new_G3453_ & new_G3431_;
  assign new_G6645_ = ~new_G6639_;
  assign new_G3470_ = ~new_G6639_ | ~new_G6646_;
  assign new_G6653_ = ~new_G6647_;
  assign new_G3473_ = ~new_G6647_ | ~new_G6654_;
  assign new_G6661_ = ~new_G6655_;
  assign new_G3477_ = ~new_G6655_ | ~new_G6662_;
  assign new_G6669_ = ~new_G6663_;
  assign new_G3480_ = ~new_G6663_ | ~new_G6670_;
  assign new_G3484_ = ~new_G6671_ | ~new_G6678_;
  assign new_G3488_ = ~new_G6679_ | ~new_G6686_;
  assign new_G3601_ = new_G3582_ & new_G3531_ & new_G3536_;
  assign new_G3604_ = new_G3586_ & new_G3527_ & new_G3540_;
  assign new_G3607_ = new_G3590_ & new_G3554_ & new_G3559_;
  assign new_G3610_ = new_G3594_ & new_G3550_ & new_G3563_;
  assign new_G4032_ = ~new_G4028_;
  assign new_G4090_ = new_G4004_ & new_G4028_;
  assign new_G4271_ = new_G4250_ & new_G4184_ & new_G4189_;
  assign new_G4274_ = new_G4254_ & new_G4180_ & new_G4193_;
  assign new_G4277_ = new_G4258_ & new_G4207_ & new_G4212_;
  assign new_G4280_ = new_G4262_ & new_G4203_ & new_G4216_;
  assign new_G4368_ = ~new_G4364_;
  assign new_G4379_ = ~new_G4376_;
  assign new_G4387_ = new_G4356_ & new_G4376_;
  assign new_G4628_ = new_G4609_ & new_G4558_ & new_G4563_;
  assign new_G4631_ = new_G4613_ & new_G4554_ & new_G4567_;
  assign new_G4634_ = new_G4617_ & new_G4581_ & new_G4586_;
  assign new_G4637_ = new_G4621_ & new_G4577_ & new_G4590_;
  assign new_G4841_ = new_G2522_ | new_G2520_ | new_G2519_ | new_G2431_ | new_G2518_;
  assign new_G4849_ = new_G2526_ | new_G2524_ | new_G2448_ | new_G2523_;
  assign new_G4857_ = new_G2529_ | new_G2465_ | new_G2527_;
  assign new_G4865_ = new_G2481_ | new_G2531_;
  assign new_G5021_ = ~new_G5019_ | ~new_G5020_;
  assign new_G5028_ = ~new_G5024_;
  assign new_G5109_ = ~new_G5107_ | ~new_G5108_;
  assign new_G5116_ = ~new_G5112_;
  assign new_G5369_ = ~new_G1313_ | ~new_G1310_;
  assign new_G5377_ = ~new_G1319_ | ~new_G1316_;
  assign new_G5385_ = ~new_G1325_ | ~new_G1322_;
  assign new_G5472_ = ~new_G5468_;
  assign new_G5473_ = ~new_G5468_ | ~new_G5471_;
  assign new_G5530_ = ~new_G5526_;
  assign new_G5531_ = ~new_G5526_ | ~new_G5529_;
  assign new_G5591_ = ~new_G5589_ | ~new_G5590_;
  assign new_G5598_ = ~new_G5594_;
  assign new_G5679_ = ~new_G5677_ | ~new_G5678_;
  assign new_G5686_ = ~new_G5682_;
  assign new_G6060_ = new_G2768_ | new_G2804_;
  assign new_G6074_ = ~new_G6070_;
  assign new_G6118_ = ~new_G2768_;
  assign new_G6132_ = ~new_G6128_;
  assign new_G6176_ = new_G2797_ | new_G2796_ | new_G2693_ | new_G2795_;
  assign new_G6186_ = new_G2801_ | new_G2807_;
  assign new_G6196_ = new_G2791_ | new_G2790_ | new_G2789_ | new_G2670_ | new_G2788_;
  assign new_G6268_ = ~new_G6264_;
  assign new_G6269_ = ~new_G6264_ | ~new_G6267_;
  assign new_G6274_ = ~new_G2801_;
  assign new_G6288_ = ~new_G6284_;
  assign new_G6337_ = ~new_G4288_ | ~new_G4285_;
  assign new_G6829_ = ~new_G3600_ | ~new_G3597_;
  assign new_G6928_ = new_G4017_ | new_G4051_;
  assign new_G6942_ = ~new_G6938_;
  assign new_G6986_ = ~new_G4017_;
  assign new_G7000_ = ~new_G6996_;
  assign new_G7048_ = ~new_G7044_;
  assign new_G7049_ = ~new_G7044_ | ~new_G7047_;
  assign new_G7054_ = new_G4048_ | new_G4052_;
  assign new_G7068_ = ~new_G7064_;
  assign new_G7136_ = ~new_G7132_;
  assign new_G7137_ = ~new_G7132_ | ~new_G7135_;
  assign new_G7142_ = ~new_G4048_;
  assign new_G7156_ = ~new_G7152_;
  assign new_G7433_ = ~new_G4627_ | ~new_G4624_;
  assign new_G242_ = new_G1982_ & new_G1146_;
  assign new_G3151_ = ~new_G3135_ | ~new_G3127_;
  assign new_G257_ = new_G3249_ & new_G3035_ & new_G3156_ & G89 & new_G4386_;
  assign new_G263_ = new_G3249_ & new_G3035_ & new_G3156_ & G89 & new_G4386_;
  assign new_G266_ = new_G1790_ & new_G997_;
  assign new_G1991_ = ~new_G1990_;
  assign new_G1998_ = ~new_G1997_;
  assign new_G3489_ = ~new_G3487_ | ~new_G3488_;
  assign new_G371_ = ~new_G4836_ | ~new_G4839_;
  assign new_G4840_ = ~new_G4836_;
  assign new_G2561_ = ~new_G2559_ | ~new_G2560_;
  assign new_G2532_ = new_G2487_ & new_G2508_;
  assign new_G2537_ = new_G2495_ | new_G2536_;
  assign new_G2541_ = ~new_G5940_ | ~new_G5943_;
  assign new_G2544_ = ~new_G5948_ | ~new_G5951_;
  assign new_G2548_ = ~new_G5956_ | ~new_G5959_;
  assign new_G2551_ = ~new_G5964_ | ~new_G5967_;
  assign new_G2557_ = ~new_G2555_ | ~new_G2556_;
  assign new_G2563_ = new_G2508_ & G4526;
  assign new_G2577_ = ~new_G2499_ | ~new_G2491_;
  assign new_G2775_ = ~new_G2771_;
  assign new_G2806_ = ~new_G2771_ | ~G4526;
  assign new_G2808_ = ~new_G2761_ | ~new_G2753_;
  assign new_G2852_ = new_G2749_ & new_G2771_;
  assign new_G2854_ = new_G2757_ | new_G2853_;
  assign new_G6366_ = ~new_G6362_;
  assign new_G4381_ = ~new_G4368_ | ~new_G4360_;
  assign new_G3164_ = new_G3131_ | new_G3163_;
  assign new_G3241_ = new_G3035_ & new_G3156_ & G89 & new_G4386_;
  assign new_G3468_ = new_G3437_ | new_G3467_;
  assign new_G3469_ = ~new_G6642_ | ~new_G6645_;
  assign new_G3472_ = ~new_G6650_ | ~new_G6653_;
  assign new_G3476_ = ~new_G6658_ | ~new_G6661_;
  assign new_G3479_ = ~new_G6666_ | ~new_G6669_;
  assign new_G3485_ = ~new_G3483_ | ~new_G3484_;
  assign new_G3603_ = ~new_G3601_ & ~new_G3602_;
  assign new_G3606_ = ~new_G3604_ & ~new_G3605_;
  assign new_G3609_ = ~new_G3607_ & ~new_G3608_;
  assign new_G3612_ = ~new_G3610_ & ~new_G3611_;
  assign new_G6844_ = ~new_G6840_;
  assign new_G6852_ = ~new_G6848_;
  assign new_G4091_ = new_G4010_ | new_G4090_;
  assign new_G4273_ = ~new_G4271_ & ~new_G4272_;
  assign new_G4276_ = ~new_G4274_ & ~new_G4275_;
  assign new_G4279_ = ~new_G4277_ & ~new_G4278_;
  assign new_G4282_ = ~new_G4280_ & ~new_G4281_;
  assign new_G4382_ = new_G4379_ & new_G4380_;
  assign new_G4388_ = new_G4364_ | new_G4387_;
  assign new_G7452_ = ~new_G7448_;
  assign new_G7462_ = ~new_G7458_;
  assign new_G4630_ = ~new_G4628_ & ~new_G4629_;
  assign new_G4633_ = ~new_G4631_ & ~new_G4632_;
  assign new_G4636_ = ~new_G4634_ & ~new_G4635_;
  assign new_G4639_ = ~new_G4637_ & ~new_G4638_;
  assign new_G4955_ = ~new_G4949_;
  assign new_G4958_ = ~new_G4949_ | ~new_G4956_;
  assign new_G4996_ = ~new_G4990_;
  assign new_G4999_ = ~new_G4990_ | ~new_G4997_;
  assign new_G5474_ = ~new_G5465_ | ~new_G5472_;
  assign new_G5532_ = ~new_G5523_ | ~new_G5530_;
  assign new_G6210_ = ~new_G6206_;
  assign new_G6270_ = ~new_G6261_ | ~new_G6268_;
  assign new_G6298_ = ~new_G6294_;
  assign new_G7050_ = ~new_G7041_ | ~new_G7048_;
  assign new_G7138_ = ~new_G7129_ | ~new_G7136_;
  assign new_G3471_ = ~new_G3469_ | ~new_G3470_;
  assign new_G3478_ = ~new_G3476_ | ~new_G3477_;
  assign new_G3486_ = ~new_G3485_;
  assign new_G372_ = ~new_G4833_ | ~new_G4840_;
  assign new_G2543_ = ~new_G2541_ | ~new_G2542_;
  assign new_G2550_ = ~new_G2548_ | ~new_G2549_;
  assign new_G2558_ = ~new_G2557_;
  assign new_G4847_ = ~new_G4841_;
  assign new_G387_ = ~new_G4841_ | ~new_G4848_;
  assign new_G4855_ = ~new_G4849_;
  assign new_G390_ = ~new_G4849_ | ~new_G4856_;
  assign new_G4863_ = ~new_G4857_;
  assign new_G393_ = ~new_G4857_ | ~new_G4864_;
  assign new_G4871_ = ~new_G4865_;
  assign new_G396_ = ~new_G4865_ | ~new_G4872_;
  assign new_G965_ = ~new_G962_;
  assign new_G5375_ = ~new_G5369_;
  assign new_G1327_ = ~new_G5369_ | ~new_G5376_;
  assign new_G5383_ = ~new_G5377_;
  assign new_G1330_ = ~new_G5377_ | ~new_G5384_;
  assign new_G5391_ = ~new_G5385_;
  assign new_G1333_ = ~new_G5385_ | ~new_G5392_;
  assign new_G1754_ = ~new_G1751_;
  assign new_G2546_ = ~new_G2544_ | ~new_G2545_;
  assign new_G2553_ = ~new_G2551_ | ~new_G2552_;
  assign new_G2564_ = new_G2515_ | new_G2563_;
  assign new_G2809_ = new_G2784_ & new_G2806_;
  assign new_G2813_ = new_G2784_ & new_G2775_;
  assign new_G6345_ = ~new_G6337_;
  assign new_G2860_ = ~new_G6337_ | ~new_G6346_;
  assign new_G3474_ = ~new_G3472_ | ~new_G3473_;
  assign new_G3481_ = ~new_G3479_ | ~new_G3480_;
  assign new_G6835_ = ~new_G6829_;
  assign new_G3614_ = ~new_G6829_ | ~new_G6836_;
  assign new_G4053_ = new_G4032_ & new_G4023_;
  assign new_G7441_ = ~new_G7433_;
  assign new_G4516_ = ~new_G7433_ | ~new_G7442_;
  assign new_G4957_ = ~new_G4952_ | ~new_G4955_;
  assign new_G4998_ = ~new_G4993_ | ~new_G4996_;
  assign new_G5027_ = ~new_G5021_;
  assign new_G5030_ = ~new_G5021_ | ~new_G5028_;
  assign new_G5115_ = ~new_G5109_;
  assign new_G5118_ = ~new_G5109_ | ~new_G5116_;
  assign new_G5475_ = ~new_G5473_ | ~new_G5474_;
  assign new_G5533_ = ~new_G5531_ | ~new_G5532_;
  assign new_G5597_ = ~new_G5591_;
  assign new_G5600_ = ~new_G5591_ | ~new_G5598_;
  assign new_G5685_ = ~new_G5679_;
  assign new_G5688_ = ~new_G5679_ | ~new_G5686_;
  assign new_G6064_ = ~new_G6060_;
  assign new_G6065_ = ~new_G6060_ | ~new_G6063_;
  assign new_G6122_ = ~new_G6118_;
  assign new_G6123_ = ~new_G6118_ | ~new_G6121_;
  assign new_G6180_ = ~new_G6176_;
  assign new_G6181_ = ~new_G6176_ | ~new_G6179_;
  assign new_G6190_ = ~new_G6186_;
  assign new_G6200_ = ~new_G6196_;
  assign new_G6271_ = ~new_G6269_ | ~new_G6270_;
  assign new_G6278_ = ~new_G6274_;
  assign new_G6347_ = ~new_G4276_ | ~new_G4273_;
  assign new_G6357_ = ~new_G4282_ | ~new_G4279_;
  assign new_G6837_ = ~new_G3606_ | ~new_G3603_;
  assign new_G6845_ = ~new_G3612_ | ~new_G3609_;
  assign new_G6932_ = ~new_G6928_;
  assign new_G6933_ = ~new_G6928_ | ~new_G6931_;
  assign new_G6990_ = ~new_G6986_;
  assign new_G6991_ = ~new_G6986_ | ~new_G6989_;
  assign new_G7051_ = ~new_G7049_ | ~new_G7050_;
  assign new_G7058_ = ~new_G7054_;
  assign new_G7139_ = ~new_G7137_ | ~new_G7138_;
  assign new_G7146_ = ~new_G7142_;
  assign new_G7443_ = ~new_G4639_ | ~new_G4636_;
  assign new_G7453_ = ~new_G4633_ | ~new_G4630_;
  assign new_G243_ = new_G1146_ & new_G3468_ & new_G1974_;
  assign new_G244_ = new_G1146_ & new_G1974_ & new_G2537_ & new_G3466_;
  assign new_G245_ = new_G1146_ & new_G1974_ & new_G3466_ & G4526 & new_G2532_;
  assign new_G255_ = new_G3249_ & new_G3164_ & new_G3035_;
  assign new_G256_ = new_G3249_ & new_G3035_ & new_G4388_ & new_G3156_;
  assign new_G261_ = new_G3249_ & new_G3164_ & new_G3035_;
  assign new_G262_ = new_G3249_ & new_G3035_ & new_G4388_ & new_G3156_;
  assign new_G267_ = new_G997_ & new_G4091_ & new_G1788_;
  assign new_G268_ = new_G997_ & new_G1788_ & new_G2854_ & new_G4089_;
  assign new_G269_ = new_G997_ & new_G1788_ & new_G4089_ & G4526 & new_G2852_;
  assign new_G3475_ = ~new_G3474_;
  assign new_G3482_ = ~new_G3481_;
  assign G373 = ~new_G371_ | ~new_G372_;
  assign new_G2547_ = ~new_G2546_;
  assign new_G2554_ = ~new_G2553_;
  assign new_G386_ = ~new_G4844_ | ~new_G4847_;
  assign new_G389_ = ~new_G4852_ | ~new_G4855_;
  assign new_G392_ = ~new_G4860_ | ~new_G4863_;
  assign new_G395_ = ~new_G4868_ | ~new_G4871_;
  assign new_G1326_ = ~new_G5372_ | ~new_G5375_;
  assign new_G1329_ = ~new_G5380_ | ~new_G5383_;
  assign new_G1332_ = ~new_G5388_ | ~new_G5391_;
  assign new_G1436_ = new_G4091_ & new_G1788_;
  assign new_G1440_ = new_G1788_ & new_G2854_ & new_G4089_;
  assign new_G1445_ = new_G1788_ & new_G4089_ & G4526 & new_G2852_;
  assign new_G1450_ = new_G2854_ & new_G4089_;
  assign new_G1454_ = new_G4089_ & G4526 & new_G2852_;
  assign new_G2859_ = ~new_G6342_ | ~new_G6345_;
  assign new_G4385_ = ~new_G4382_;
  assign new_G3148_ = new_G4382_ & new_G4364_;
  assign new_G3239_ = new_G3164_ & new_G3035_;
  assign new_G3240_ = new_G3035_ & new_G4388_ & new_G3156_;
  assign new_G3265_ = new_G3468_ & new_G1974_;
  assign new_G3267_ = new_G1974_ & new_G2537_ & new_G3466_;
  assign new_G3270_ = new_G1974_ & new_G3466_ & G4526 & new_G2532_;
  assign new_G3274_ = new_G2537_ & new_G3466_;
  assign new_G3277_ = new_G3466_ & G4526 & new_G2532_;
  assign new_G3613_ = ~new_G6832_ | ~new_G6835_;
  assign new_G4515_ = ~new_G7438_ | ~new_G7441_;
  assign new_G4959_ = ~new_G4957_ | ~new_G4958_;
  assign new_G5000_ = ~new_G4998_ | ~new_G4999_;
  assign new_G5029_ = ~new_G5024_ | ~new_G5027_;
  assign new_G5117_ = ~new_G5112_ | ~new_G5115_;
  assign new_G5599_ = ~new_G5594_ | ~new_G5597_;
  assign new_G5687_ = ~new_G5682_ | ~new_G5685_;
  assign new_G6066_ = ~new_G6057_ | ~new_G6064_;
  assign new_G6124_ = ~new_G6115_ | ~new_G6122_;
  assign new_G6182_ = ~new_G6173_ | ~new_G6180_;
  assign new_G6934_ = ~new_G6925_ | ~new_G6932_;
  assign new_G6992_ = ~new_G6983_ | ~new_G6990_;
  assign G246 = new_G245_ | new_G244_ | new_G243_ | new_G241_ | new_G242_;
  assign G258 = new_G257_ | new_G256_ | new_G255_ | new_G3259_ | new_G254_;
  assign G264 = new_G263_ | new_G262_ | new_G261_ | new_G3259_ | new_G260_;
  assign G270 = new_G269_ | new_G268_ | new_G267_ | new_G265_ | new_G266_;
  assign new_G375_ = new_G2564_ & new_G2543_;
  assign new_G378_ = new_G2564_ & new_G2550_;
  assign new_G381_ = new_G2564_ & new_G2558_;
  assign new_G384_ = new_G2564_ & new_G2406_;
  assign G388 = ~new_G386_ | ~new_G387_;
  assign G391 = ~new_G389_ | ~new_G390_;
  assign G394 = ~new_G392_ | ~new_G393_;
  assign G397 = ~new_G395_ | ~new_G396_;
  assign new_G1328_ = ~new_G1326_ | ~new_G1327_;
  assign new_G1331_ = ~new_G1329_ | ~new_G1330_;
  assign new_G1334_ = ~new_G1332_ | ~new_G1333_;
  assign new_G1447_ = new_G1445_ | new_G1440_ | new_G1790_ | new_G1436_;
  assign new_G1766_ = new_G1454_ | new_G4091_ | new_G1450_;
  assign new_G2571_ = ~new_G2564_;
  assign new_G2579_ = new_G2577_ & new_G2564_;
  assign new_G2812_ = ~new_G2809_;
  assign new_G2816_ = ~new_G2813_;
  assign new_G2851_ = new_G2809_ & new_G2757_;
  assign new_G2861_ = ~new_G2859_ | ~new_G2860_;
  assign new_G6355_ = ~new_G6347_;
  assign new_G2863_ = ~new_G6347_ | ~new_G6356_;
  assign new_G6365_ = ~new_G6357_;
  assign new_G2866_ = ~new_G6357_ | ~new_G6366_;
  assign new_G3147_ = new_G4381_ & new_G4385_;
  assign new_G3242_ = new_G3241_ | new_G3240_ | new_G3046_ | new_G3239_;
  assign new_G3271_ = new_G3270_ | new_G3267_ | new_G1982_ | new_G3265_;
  assign new_G3279_ = new_G3277_ | new_G3468_ | new_G3274_;
  assign new_G3615_ = ~new_G3613_ | ~new_G3614_;
  assign new_G6843_ = ~new_G6837_;
  assign new_G3617_ = ~new_G6837_ | ~new_G6844_;
  assign new_G6851_ = ~new_G6845_;
  assign new_G3620_ = ~new_G6845_ | ~new_G6852_;
  assign new_G4056_ = ~new_G4053_;
  assign new_G4517_ = ~new_G4515_ | ~new_G4516_;
  assign new_G7451_ = ~new_G7443_;
  assign new_G4519_ = ~new_G7443_ | ~new_G7452_;
  assign new_G7461_ = ~new_G7453_;
  assign new_G4522_ = ~new_G7453_ | ~new_G7462_;
  assign new_G5031_ = ~new_G5029_ | ~new_G5030_;
  assign new_G5119_ = ~new_G5117_ | ~new_G5118_;
  assign new_G5481_ = ~new_G5475_;
  assign new_G5484_ = ~new_G5475_ | ~new_G5482_;
  assign new_G5539_ = ~new_G5533_;
  assign new_G5542_ = ~new_G5533_ | ~new_G5540_;
  assign new_G5601_ = ~new_G5599_ | ~new_G5600_;
  assign new_G5689_ = ~new_G5687_ | ~new_G5688_;
  assign new_G6067_ = ~new_G6065_ | ~new_G6066_;
  assign new_G6125_ = ~new_G6123_ | ~new_G6124_;
  assign new_G6183_ = ~new_G6181_ | ~new_G6182_;
  assign new_G6277_ = ~new_G6271_;
  assign new_G6280_ = ~new_G6271_ | ~new_G6278_;
  assign new_G6935_ = ~new_G6933_ | ~new_G6934_;
  assign new_G6993_ = ~new_G6991_ | ~new_G6992_;
  assign new_G7057_ = ~new_G7051_;
  assign new_G7060_ = ~new_G7051_ | ~new_G7058_;
  assign new_G7145_ = ~new_G7139_;
  assign new_G7148_ = ~new_G7139_ | ~new_G7146_;
  assign new_G4968_ = ~new_G4959_ | ~new_G4966_;
  assign new_G5009_ = ~new_G5000_ | ~new_G5007_;
  assign new_G2850_ = new_G2808_ & new_G2812_;
  assign new_G2862_ = ~new_G6352_ | ~new_G6355_;
  assign new_G2865_ = ~new_G6362_ | ~new_G6365_;
  assign new_G3149_ = new_G3147_ | new_G3148_;
  assign new_G3243_ = ~new_G3228_ | ~new_G3242_;
  assign new_G3616_ = ~new_G6840_ | ~new_G6843_;
  assign new_G3619_ = ~new_G6848_ | ~new_G6851_;
  assign new_G4518_ = ~new_G7448_ | ~new_G7451_;
  assign new_G4521_ = ~new_G7458_ | ~new_G7461_;
  assign new_G4965_ = ~new_G4959_;
  assign new_G5006_ = ~new_G5000_;
  assign new_G5483_ = ~new_G5478_ | ~new_G5481_;
  assign new_G5541_ = ~new_G5536_ | ~new_G5539_;
  assign new_G6279_ = ~new_G6274_ | ~new_G6277_;
  assign new_G7059_ = ~new_G7054_ | ~new_G7057_;
  assign new_G7147_ = ~new_G7142_ | ~new_G7145_;
  assign new_G374_ = new_G2547_ & new_G2571_;
  assign new_G377_ = new_G2554_ & new_G2571_;
  assign new_G380_ = new_G2561_ & new_G2571_;
  assign new_G383_ = new_G2400_ & new_G2571_;
  assign new_G955_ = ~new_G920_ | ~new_G1447_;
  assign new_G4967_ = ~new_G4962_ | ~new_G4965_;
  assign new_G5008_ = ~new_G5003_ | ~new_G5006_;
  assign new_G975_ = new_G1447_;
  assign new_G1136_ = new_G1038_ & new_G1074_ & new_G1055_ & new_G3271_ & new_G1093_;
  assign new_G1140_ = new_G1074_ & new_G1055_ & new_G3271_ & new_G1093_;
  assign new_G1143_ = new_G1074_ & new_G3271_ & new_G1093_;
  assign new_G1145_ = new_G3271_ & new_G1093_;
  assign new_G1160_ = new_G1122_ & new_G3271_;
  assign new_G1771_ = ~new_G1766_;
  assign new_G1964_ = new_G1869_ & new_G1903_ & new_G1885_ & new_G3279_ & new_G1921_;
  assign new_G1968_ = new_G1903_ & new_G1885_ & new_G3279_ & new_G1921_;
  assign new_G1971_ = new_G1903_ & new_G3279_ & new_G1921_;
  assign new_G1973_ = new_G3279_ & new_G1921_;
  assign new_G2007_ = new_G1950_ & new_G3279_;
  assign new_G2578_ = new_G2495_ & new_G2571_;
  assign new_G2864_ = ~new_G2862_ | ~new_G2863_;
  assign new_G2867_ = ~new_G2865_ | ~new_G2866_;
  assign new_G3150_ = ~new_G3136_ | ~new_G3149_;
  assign new_G3245_ = new_G3238_ & new_G3243_;
  assign new_G3618_ = ~new_G3616_ | ~new_G3617_;
  assign new_G3621_ = ~new_G3619_ | ~new_G3620_;
  assign new_G4067_ = new_G2850_ | new_G2851_;
  assign new_G4520_ = ~new_G4518_ | ~new_G4519_;
  assign new_G4523_ = ~new_G4521_ | ~new_G4522_;
  assign new_G4713_ = new_G3279_;
  assign new_G4753_ = new_G3271_;
  assign new_G5037_ = ~new_G5031_;
  assign new_G5040_ = ~new_G5031_ | ~new_G5038_;
  assign new_G5125_ = ~new_G5119_;
  assign new_G5128_ = ~new_G5119_ | ~new_G5126_;
  assign new_G5485_ = ~new_G5483_ | ~new_G5484_;
  assign new_G5543_ = ~new_G5541_ | ~new_G5542_;
  assign new_G5607_ = ~new_G5601_;
  assign new_G5610_ = ~new_G5601_ | ~new_G5608_;
  assign new_G5695_ = ~new_G5689_;
  assign new_G5698_ = ~new_G5689_ | ~new_G5696_;
  assign new_G6073_ = ~new_G6067_;
  assign new_G6076_ = ~new_G6067_ | ~new_G6074_;
  assign new_G6131_ = ~new_G6125_;
  assign new_G6134_ = ~new_G6125_ | ~new_G6132_;
  assign new_G6189_ = ~new_G6183_;
  assign new_G6192_ = ~new_G6183_ | ~new_G6190_;
  assign new_G6281_ = ~new_G6279_ | ~new_G6280_;
  assign new_G6941_ = ~new_G6935_;
  assign new_G6944_ = ~new_G6935_ | ~new_G6942_;
  assign new_G6999_ = ~new_G6993_;
  assign new_G7002_ = ~new_G6993_ | ~new_G7000_;
  assign new_G7061_ = ~new_G7059_ | ~new_G7060_;
  assign new_G7149_ = ~new_G7147_ | ~new_G7148_;
  assign G376 = new_G374_ | new_G375_;
  assign G379 = new_G377_ | new_G378_;
  assign G382 = new_G380_ | new_G381_;
  assign G385 = new_G383_ | new_G384_;
  assign new_G958_ = new_G933_ & new_G955_;
  assign new_G967_ = ~new_G4967_ | ~new_G4968_;
  assign new_G971_ = ~new_G5008_ | ~new_G5009_;
  assign new_G1161_ = new_G1129_ | new_G1160_;
  assign new_G2008_ = new_G1957_ | new_G2007_;
  assign new_G2580_ = new_G2578_ | new_G2579_;
  assign new_G2868_ = new_G2867_ & new_G2864_ & new_G1331_ & new_G2861_;
  assign new_G3152_ = new_G3146_ & new_G3150_;
  assign new_G4443_ = new_G3621_ & new_G3618_ & new_G1328_ & new_G1334_;
  assign new_G4524_ = new_G4523_ & new_G4520_ & new_G3615_ & new_G4517_;
  assign new_G4721_ = new_G1964_ | new_G1962_ | new_G1961_ | new_G1880_ | new_G1960_;
  assign new_G4729_ = new_G1968_ | new_G1966_ | new_G1897_ | new_G1965_;
  assign new_G4737_ = new_G1971_ | new_G1914_ | new_G1969_;
  assign new_G4745_ = new_G1929_ | new_G1973_;
  assign new_G4761_ = new_G1136_ | new_G1134_ | new_G1133_ | new_G1050_ | new_G1132_;
  assign new_G4769_ = new_G1140_ | new_G1138_ | new_G1068_ | new_G1137_;
  assign new_G4777_ = new_G1143_ | new_G1086_ | new_G1141_;
  assign new_G4785_ = new_G1102_ | new_G1145_;
  assign new_G5039_ = ~new_G5034_ | ~new_G5037_;
  assign new_G5127_ = ~new_G5122_ | ~new_G5125_;
  assign new_G5609_ = ~new_G5604_ | ~new_G5607_;
  assign new_G5697_ = ~new_G5692_ | ~new_G5695_;
  assign new_G6075_ = ~new_G6070_ | ~new_G6073_;
  assign new_G6133_ = ~new_G6128_ | ~new_G6131_;
  assign new_G6191_ = ~new_G6186_ | ~new_G6189_;
  assign new_G6943_ = ~new_G6938_ | ~new_G6941_;
  assign new_G7001_ = ~new_G6996_ | ~new_G6999_;
  assign new_G3248_ = ~new_G3245_;
  assign new_G248_ = new_G3245_ & new_G3223_;
  assign new_G4719_ = ~new_G4713_;
  assign new_G294_ = ~new_G4713_ | ~new_G4720_;
  assign new_G4759_ = ~new_G4753_;
  assign new_G323_ = ~new_G4753_ | ~new_G4760_;
  assign new_G980_ = ~new_G975_;
  assign new_G4072_ = ~new_G4067_;
  assign new_G5041_ = ~new_G5039_ | ~new_G5040_;
  assign new_G5129_ = ~new_G5127_ | ~new_G5128_;
  assign new_G5491_ = ~new_G5485_;
  assign new_G5494_ = ~new_G5485_ | ~new_G5492_;
  assign new_G5549_ = ~new_G5543_;
  assign new_G5552_ = ~new_G5543_ | ~new_G5550_;
  assign new_G5611_ = ~new_G5609_ | ~new_G5610_;
  assign new_G5699_ = ~new_G5697_ | ~new_G5698_;
  assign new_G6077_ = ~new_G6075_ | ~new_G6076_;
  assign new_G6135_ = ~new_G6133_ | ~new_G6134_;
  assign new_G6193_ = ~new_G6191_ | ~new_G6192_;
  assign new_G6287_ = ~new_G6281_;
  assign new_G6290_ = ~new_G6281_ | ~new_G6288_;
  assign new_G6945_ = ~new_G6943_ | ~new_G6944_;
  assign new_G7003_ = ~new_G7001_ | ~new_G7002_;
  assign new_G7067_ = ~new_G7061_;
  assign new_G7070_ = ~new_G7061_ | ~new_G7068_;
  assign new_G7155_ = ~new_G7149_;
  assign new_G7158_ = ~new_G7149_ | ~new_G7156_;
  assign new_G247_ = new_G3244_ & new_G3248_;
  assign new_G3155_ = ~new_G3152_;
  assign new_G251_ = new_G3152_ & new_G3131_;
  assign new_G272_ = new_G1176_ & new_G1161_;
  assign new_G961_ = ~new_G958_;
  assign new_G275_ = new_G958_ & new_G908_;
  assign new_G293_ = ~new_G4716_ | ~new_G4719_;
  assign new_G297_ = new_G2008_ & new_G1987_;
  assign new_G300_ = new_G2008_ & new_G1994_;
  assign new_G303_ = new_G2008_ & new_G2002_;
  assign new_G306_ = new_G2008_ & new_G1856_;
  assign new_G4727_ = ~new_G4721_;
  assign new_G309_ = ~new_G4721_ | ~new_G4728_;
  assign new_G4735_ = ~new_G4729_;
  assign new_G312_ = ~new_G4729_ | ~new_G4736_;
  assign new_G4743_ = ~new_G4737_;
  assign new_G315_ = ~new_G4737_ | ~new_G4744_;
  assign new_G4751_ = ~new_G4745_;
  assign new_G318_ = ~new_G4745_ | ~new_G4752_;
  assign new_G322_ = ~new_G4756_ | ~new_G4759_;
  assign new_G4767_ = ~new_G4761_;
  assign new_G326_ = ~new_G4761_ | ~new_G4768_;
  assign new_G4775_ = ~new_G4769_;
  assign new_G329_ = ~new_G4769_ | ~new_G4776_;
  assign new_G4783_ = ~new_G4777_;
  assign new_G332_ = ~new_G4777_ | ~new_G4784_;
  assign new_G4791_ = ~new_G4785_;
  assign new_G335_ = ~new_G4785_ | ~new_G4792_;
  assign G412 = ~new_G4443_;
  assign G414 = ~new_G4524_;
  assign G416 = ~new_G2868_;
  assign new_G2881_ = new_G2868_ & new_G4443_ & new_G4524_;
  assign new_G993_ = new_G975_ & new_G971_ & new_G962_;
  assign new_G994_ = new_G975_ & new_G967_ & new_G965_;
  assign new_G1166_ = ~new_G1161_;
  assign new_G1171_ = new_G1161_ & new_G1155_;
  assign new_G1174_ = new_G1161_ & new_G1023_;
  assign new_G2014_ = ~new_G2008_;
  assign new_G3459_ = new_G3365_ & new_G3399_ & new_G3381_ & new_G2580_ & new_G3417_;
  assign new_G3462_ = new_G3399_ & new_G3381_ & new_G2580_ & new_G3417_;
  assign new_G3464_ = new_G3399_ & new_G2580_ & new_G3417_;
  assign new_G3465_ = new_G2580_ & new_G3417_;
  assign new_G3490_ = new_G3446_ & new_G2580_;
  assign new_G4793_ = new_G2580_;
  assign new_G5493_ = ~new_G5488_ | ~new_G5491_;
  assign new_G5551_ = ~new_G5546_ | ~new_G5549_;
  assign new_G6289_ = ~new_G6284_ | ~new_G6287_;
  assign new_G7069_ = ~new_G7064_ | ~new_G7067_;
  assign new_G7157_ = ~new_G7152_ | ~new_G7155_;
  assign G249 = new_G247_ | new_G248_;
  assign new_G250_ = new_G3151_ & new_G3155_;
  assign new_G274_ = new_G957_ & new_G961_;
  assign G295 = ~new_G293_ | ~new_G294_;
  assign new_G308_ = ~new_G4724_ | ~new_G4727_;
  assign new_G311_ = ~new_G4732_ | ~new_G4735_;
  assign new_G314_ = ~new_G4740_ | ~new_G4743_;
  assign new_G317_ = ~new_G4748_ | ~new_G4751_;
  assign G324 = ~new_G322_ | ~new_G323_;
  assign new_G325_ = ~new_G4764_ | ~new_G4767_;
  assign new_G328_ = ~new_G4772_ | ~new_G4775_;
  assign new_G331_ = ~new_G4780_ | ~new_G4783_;
  assign new_G334_ = ~new_G4788_ | ~new_G4791_;
  assign new_G417_ = new_G2881_ & new_G2876_ & new_G2878_;
  assign new_G991_ = new_G980_ & new_G971_ & new_G933_;
  assign new_G992_ = new_G980_ & new_G967_ & new_G929_;
  assign new_G3491_ = new_G3453_ | new_G3490_;
  assign new_G4801_ = new_G3459_ | new_G3458_ | new_G3457_ | new_G3376_ | new_G3456_;
  assign new_G4809_ = new_G3462_ | new_G3461_ | new_G3393_ | new_G3460_;
  assign new_G4817_ = new_G3464_ | new_G3410_ | new_G3463_;
  assign new_G4825_ = new_G3425_ | new_G3465_;
  assign new_G5047_ = ~new_G5041_;
  assign new_G5050_ = ~new_G5041_ | ~new_G5048_;
  assign new_G5135_ = ~new_G5129_;
  assign new_G5138_ = ~new_G5129_ | ~new_G5136_;
  assign new_G5495_ = ~new_G5493_ | ~new_G5494_;
  assign new_G5553_ = ~new_G5551_ | ~new_G5552_;
  assign new_G5617_ = ~new_G5611_;
  assign new_G5620_ = ~new_G5611_ | ~new_G5618_;
  assign new_G5705_ = ~new_G5699_;
  assign new_G5708_ = ~new_G5699_ | ~new_G5706_;
  assign new_G6083_ = ~new_G6077_;
  assign new_G6086_ = ~new_G6077_ | ~new_G6084_;
  assign new_G6141_ = ~new_G6135_;
  assign new_G6144_ = ~new_G6135_ | ~new_G6142_;
  assign new_G6199_ = ~new_G6193_;
  assign new_G6202_ = ~new_G6193_ | ~new_G6200_;
  assign new_G6291_ = ~new_G6289_ | ~new_G6290_;
  assign new_G6951_ = ~new_G6945_;
  assign new_G6954_ = ~new_G6945_ | ~new_G6952_;
  assign new_G7009_ = ~new_G7003_;
  assign new_G7012_ = ~new_G7003_ | ~new_G7010_;
  assign new_G7071_ = ~new_G7069_ | ~new_G7070_;
  assign new_G7159_ = ~new_G7157_ | ~new_G7158_;
  assign G252 = new_G250_ | new_G251_;
  assign new_G271_ = new_G1117_ & new_G1166_;
  assign G276 = new_G274_ | new_G275_;
  assign new_G296_ = new_G1991_ & new_G2014_;
  assign new_G299_ = new_G1998_ & new_G2014_;
  assign new_G302_ = new_G2005_ & new_G2014_;
  assign new_G305_ = new_G1850_ & new_G2014_;
  assign G310 = ~new_G308_ | ~new_G309_;
  assign G313 = ~new_G311_ | ~new_G312_;
  assign G316 = ~new_G314_ | ~new_G315_;
  assign G319 = ~new_G317_ | ~new_G318_;
  assign G327 = ~new_G325_ | ~new_G326_;
  assign G330 = ~new_G328_ | ~new_G329_;
  assign G333 = ~new_G331_ | ~new_G332_;
  assign G336 = ~new_G334_ | ~new_G335_;
  assign new_G4799_ = ~new_G4793_;
  assign new_G343_ = ~new_G4793_ | ~new_G4800_;
  assign G418 = ~new_G417_;
  assign new_G1170_ = new_G1158_ & new_G1166_;
  assign new_G1173_ = new_G1019_ & new_G1166_;
  assign new_G5049_ = ~new_G5044_ | ~new_G5047_;
  assign new_G5137_ = ~new_G5132_ | ~new_G5135_;
  assign new_G5167_ = new_G994_ | new_G993_ | new_G991_ | new_G992_;
  assign new_G5619_ = ~new_G5614_ | ~new_G5617_;
  assign new_G5707_ = ~new_G5702_ | ~new_G5705_;
  assign new_G6085_ = ~new_G6080_ | ~new_G6083_;
  assign new_G6143_ = ~new_G6138_ | ~new_G6141_;
  assign new_G6201_ = ~new_G6196_ | ~new_G6199_;
  assign new_G6953_ = ~new_G6948_ | ~new_G6951_;
  assign new_G7011_ = ~new_G7006_ | ~new_G7009_;
  assign G273 = new_G271_ | new_G272_;
  assign G298 = new_G296_ | new_G297_;
  assign G301 = new_G299_ | new_G300_;
  assign G304 = new_G302_ | new_G303_;
  assign G307 = new_G305_ | new_G306_;
  assign new_G342_ = ~new_G4796_ | ~new_G4799_;
  assign new_G346_ = new_G3491_ & new_G3471_;
  assign new_G349_ = new_G3491_ & new_G3478_;
  assign new_G352_ = new_G3491_ & new_G3486_;
  assign new_G355_ = new_G3491_ & new_G3350_;
  assign new_G4807_ = ~new_G4801_;
  assign new_G358_ = ~new_G4801_ | ~new_G4808_;
  assign new_G4815_ = ~new_G4809_;
  assign new_G361_ = ~new_G4809_ | ~new_G4816_;
  assign new_G4823_ = ~new_G4817_;
  assign new_G364_ = ~new_G4817_ | ~new_G4824_;
  assign new_G4831_ = ~new_G4825_;
  assign new_G367_ = ~new_G4825_ | ~new_G4832_;
  assign new_G1172_ = new_G1170_ | new_G1171_;
  assign new_G1175_ = new_G1173_ | new_G1174_;
  assign new_G3497_ = ~new_G3491_;
  assign new_G5051_ = ~new_G5049_ | ~new_G5050_;
  assign new_G5139_ = ~new_G5137_ | ~new_G5138_;
  assign new_G5501_ = ~new_G5495_;
  assign new_G5504_ = ~new_G5495_ | ~new_G5502_;
  assign new_G5559_ = ~new_G5553_;
  assign new_G5562_ = ~new_G5553_ | ~new_G5560_;
  assign new_G5621_ = ~new_G5619_ | ~new_G5620_;
  assign new_G5709_ = ~new_G5707_ | ~new_G5708_;
  assign new_G6087_ = ~new_G6085_ | ~new_G6086_;
  assign new_G6145_ = ~new_G6143_ | ~new_G6144_;
  assign new_G6203_ = ~new_G6201_ | ~new_G6202_;
  assign new_G6297_ = ~new_G6291_;
  assign new_G6300_ = ~new_G6291_ | ~new_G6298_;
  assign new_G6955_ = ~new_G6953_ | ~new_G6954_;
  assign new_G7013_ = ~new_G7011_ | ~new_G7012_;
  assign new_G7077_ = ~new_G7071_;
  assign new_G7080_ = ~new_G7071_ | ~new_G7078_;
  assign new_G7165_ = ~new_G7159_;
  assign new_G7168_ = ~new_G7159_ | ~new_G7166_;
  assign G344 = ~new_G342_ | ~new_G343_;
  assign new_G357_ = ~new_G4804_ | ~new_G4807_;
  assign new_G360_ = ~new_G4812_ | ~new_G4815_;
  assign new_G363_ = ~new_G4820_ | ~new_G4823_;
  assign new_G366_ = ~new_G4828_ | ~new_G4831_;
  assign new_G5173_ = ~new_G5167_;
  assign G422 = new_G1172_;
  assign G469 = new_G1172_;
  assign G419 = new_G1175_;
  assign G471 = new_G1175_;
  assign new_G5503_ = ~new_G5498_ | ~new_G5501_;
  assign new_G5561_ = ~new_G5556_ | ~new_G5559_;
  assign new_G6299_ = ~new_G6294_ | ~new_G6297_;
  assign new_G7079_ = ~new_G7074_ | ~new_G7077_;
  assign new_G7167_ = ~new_G7162_ | ~new_G7165_;
  assign new_G345_ = new_G3475_ & new_G3497_;
  assign new_G348_ = new_G3482_ & new_G3497_;
  assign new_G351_ = new_G3489_ & new_G3497_;
  assign new_G354_ = new_G3344_ & new_G3497_;
  assign G359 = ~new_G357_ | ~new_G358_;
  assign G362 = ~new_G360_ | ~new_G361_;
  assign G365 = ~new_G363_ | ~new_G364_;
  assign G368 = ~new_G366_ | ~new_G367_;
  assign new_G5057_ = ~new_G5051_;
  assign new_G5060_ = ~new_G5051_ | ~new_G5058_;
  assign new_G5145_ = ~new_G5139_;
  assign new_G5148_ = ~new_G5139_ | ~new_G5146_;
  assign new_G5505_ = ~new_G5503_ | ~new_G5504_;
  assign new_G5563_ = ~new_G5561_ | ~new_G5562_;
  assign new_G5627_ = ~new_G5621_;
  assign new_G5630_ = ~new_G5621_ | ~new_G5628_;
  assign new_G5715_ = ~new_G5709_;
  assign new_G5718_ = ~new_G5709_ | ~new_G5716_;
  assign new_G6093_ = ~new_G6087_;
  assign new_G6096_ = ~new_G6087_ | ~new_G6094_;
  assign new_G6151_ = ~new_G6145_;
  assign new_G6154_ = ~new_G6145_ | ~new_G6152_;
  assign new_G6209_ = ~new_G6203_;
  assign new_G6212_ = ~new_G6203_ | ~new_G6210_;
  assign new_G6301_ = ~new_G6299_ | ~new_G6300_;
  assign new_G6961_ = ~new_G6955_;
  assign new_G6964_ = ~new_G6955_ | ~new_G6962_;
  assign new_G7019_ = ~new_G7013_;
  assign new_G7022_ = ~new_G7013_ | ~new_G7020_;
  assign new_G7081_ = ~new_G7079_ | ~new_G7080_;
  assign new_G7169_ = ~new_G7167_ | ~new_G7168_;
  assign G347 = new_G345_ | new_G346_;
  assign G350 = new_G348_ | new_G349_;
  assign G353 = new_G351_ | new_G352_;
  assign G356 = new_G354_ | new_G355_;
  assign new_G5059_ = ~new_G5054_ | ~new_G5057_;
  assign new_G5147_ = ~new_G5142_ | ~new_G5145_;
  assign new_G5629_ = ~new_G5624_ | ~new_G5627_;
  assign new_G5717_ = ~new_G5712_ | ~new_G5715_;
  assign new_G6095_ = ~new_G6090_ | ~new_G6093_;
  assign new_G6153_ = ~new_G6148_ | ~new_G6151_;
  assign new_G6211_ = ~new_G6206_ | ~new_G6209_;
  assign new_G6963_ = ~new_G6958_ | ~new_G6961_;
  assign new_G7021_ = ~new_G7016_ | ~new_G7019_;
  assign new_G5061_ = ~new_G5059_ | ~new_G5060_;
  assign new_G5149_ = ~new_G5147_ | ~new_G5148_;
  assign new_G5511_ = ~new_G5505_;
  assign new_G5514_ = ~new_G5505_ | ~new_G5512_;
  assign new_G5569_ = ~new_G5563_;
  assign new_G5572_ = ~new_G5563_ | ~new_G5570_;
  assign new_G5631_ = ~new_G5629_ | ~new_G5630_;
  assign new_G5719_ = ~new_G5717_ | ~new_G5718_;
  assign new_G6097_ = ~new_G6095_ | ~new_G6096_;
  assign new_G6155_ = ~new_G6153_ | ~new_G6154_;
  assign new_G6213_ = ~new_G6211_ | ~new_G6212_;
  assign new_G6307_ = ~new_G6301_;
  assign new_G6310_ = ~new_G6301_ | ~new_G6308_;
  assign new_G6965_ = ~new_G6963_ | ~new_G6964_;
  assign new_G7023_ = ~new_G7021_ | ~new_G7022_;
  assign new_G7087_ = ~new_G7081_;
  assign new_G7090_ = ~new_G7081_ | ~new_G7088_;
  assign new_G7175_ = ~new_G7169_;
  assign new_G7178_ = ~new_G7169_ | ~new_G7176_;
  assign new_G5513_ = ~new_G5508_ | ~new_G5511_;
  assign new_G5571_ = ~new_G5566_ | ~new_G5569_;
  assign new_G6309_ = ~new_G6304_ | ~new_G6307_;
  assign new_G7089_ = ~new_G7084_ | ~new_G7087_;
  assign new_G7177_ = ~new_G7172_ | ~new_G7175_;
  assign new_G5067_ = ~new_G5061_;
  assign new_G5070_ = ~new_G5061_ | ~new_G5068_;
  assign new_G5155_ = ~new_G5149_;
  assign new_G5158_ = ~new_G5149_ | ~new_G5156_;
  assign new_G5515_ = ~new_G5513_ | ~new_G5514_;
  assign new_G5573_ = ~new_G5571_ | ~new_G5572_;
  assign new_G5637_ = ~new_G5631_;
  assign new_G5640_ = ~new_G5631_ | ~new_G5638_;
  assign new_G5725_ = ~new_G5719_;
  assign new_G5728_ = ~new_G5719_ | ~new_G5726_;
  assign new_G6103_ = ~new_G6097_;
  assign new_G6106_ = ~new_G6097_ | ~new_G6104_;
  assign new_G6161_ = ~new_G6155_;
  assign new_G6164_ = ~new_G6155_ | ~new_G6162_;
  assign new_G6219_ = ~new_G6213_;
  assign new_G6222_ = ~new_G6213_ | ~new_G6220_;
  assign new_G6311_ = ~new_G6309_ | ~new_G6310_;
  assign new_G6971_ = ~new_G6965_;
  assign new_G6974_ = ~new_G6965_ | ~new_G6972_;
  assign new_G7029_ = ~new_G7023_;
  assign new_G7032_ = ~new_G7023_ | ~new_G7030_;
  assign new_G7091_ = ~new_G7089_ | ~new_G7090_;
  assign new_G7179_ = ~new_G7177_ | ~new_G7178_;
  assign new_G5069_ = ~new_G5064_ | ~new_G5067_;
  assign new_G5157_ = ~new_G5152_ | ~new_G5155_;
  assign new_G5639_ = ~new_G5634_ | ~new_G5637_;
  assign new_G5727_ = ~new_G5722_ | ~new_G5725_;
  assign new_G6105_ = ~new_G6100_ | ~new_G6103_;
  assign new_G6163_ = ~new_G6158_ | ~new_G6161_;
  assign new_G6221_ = ~new_G6216_ | ~new_G6219_;
  assign new_G6973_ = ~new_G6968_ | ~new_G6971_;
  assign new_G7031_ = ~new_G7026_ | ~new_G7029_;
  assign new_G5521_ = ~new_G5515_;
  assign new_G1756_ = ~new_G5515_ | ~new_G5522_;
  assign new_G5579_ = ~new_G5573_;
  assign new_G1761_ = ~new_G5573_ | ~new_G5580_;
  assign new_G5071_ = ~new_G5069_ | ~new_G5070_;
  assign new_G5159_ = ~new_G5157_ | ~new_G5158_;
  assign new_G5641_ = ~new_G5639_ | ~new_G5640_;
  assign new_G5729_ = ~new_G5727_ | ~new_G5728_;
  assign new_G6107_ = ~new_G6105_ | ~new_G6106_;
  assign new_G6165_ = ~new_G6163_ | ~new_G6164_;
  assign new_G6223_ = ~new_G6221_ | ~new_G6222_;
  assign new_G6317_ = ~new_G6311_;
  assign new_G6320_ = ~new_G6311_ | ~new_G6318_;
  assign new_G6975_ = ~new_G6973_ | ~new_G6974_;
  assign new_G7033_ = ~new_G7031_ | ~new_G7032_;
  assign new_G7097_ = ~new_G7091_;
  assign new_G7100_ = ~new_G7091_ | ~new_G7098_;
  assign new_G7185_ = ~new_G7179_;
  assign new_G7188_ = ~new_G7179_ | ~new_G7186_;
  assign new_G1755_ = ~new_G5518_ | ~new_G5521_;
  assign new_G1760_ = ~new_G5576_ | ~new_G5579_;
  assign new_G6319_ = ~new_G6314_ | ~new_G6317_;
  assign new_G7099_ = ~new_G7094_ | ~new_G7097_;
  assign new_G7187_ = ~new_G7182_ | ~new_G7185_;
  assign new_G1757_ = ~new_G1755_ | ~new_G1756_;
  assign new_G1762_ = ~new_G1760_ | ~new_G1761_;
  assign new_G6113_ = ~new_G6107_;
  assign new_G2818_ = ~new_G6107_ | ~new_G6114_;
  assign new_G6171_ = ~new_G6165_;
  assign new_G2823_ = ~new_G6165_ | ~new_G6172_;
  assign new_G6981_ = ~new_G6975_;
  assign new_G4058_ = ~new_G6975_ | ~new_G6982_;
  assign new_G7039_ = ~new_G7033_;
  assign new_G4063_ = ~new_G7033_ | ~new_G7040_;
  assign new_G5077_ = ~new_G5071_;
  assign new_G5080_ = ~new_G5071_ | ~new_G5078_;
  assign new_G5165_ = ~new_G5159_;
  assign new_G5090_ = ~new_G5159_ | ~new_G5166_;
  assign new_G5647_ = ~new_G5641_;
  assign new_G5650_ = ~new_G5641_ | ~new_G5648_;
  assign new_G5735_ = ~new_G5729_;
  assign new_G5660_ = ~new_G5729_ | ~new_G5736_;
  assign new_G6229_ = ~new_G6223_;
  assign new_G6232_ = ~new_G6223_ | ~new_G6230_;
  assign new_G6321_ = ~new_G6319_ | ~new_G6320_;
  assign new_G7101_ = ~new_G7099_ | ~new_G7100_;
  assign new_G7189_ = ~new_G7187_ | ~new_G7188_;
  assign new_G2817_ = ~new_G6110_ | ~new_G6113_;
  assign new_G2822_ = ~new_G6168_ | ~new_G6171_;
  assign new_G4057_ = ~new_G6978_ | ~new_G6981_;
  assign new_G4062_ = ~new_G7036_ | ~new_G7039_;
  assign new_G5079_ = ~new_G5074_ | ~new_G5077_;
  assign new_G5089_ = ~new_G5162_ | ~new_G5165_;
  assign new_G5649_ = ~new_G5644_ | ~new_G5647_;
  assign new_G5659_ = ~new_G5732_ | ~new_G5735_;
  assign new_G6231_ = ~new_G6226_ | ~new_G6229_;
  assign new_G1782_ = new_G1771_ & new_G1762_ & new_G1730_;
  assign new_G1783_ = new_G1771_ & new_G1757_ & new_G1726_;
  assign new_G1784_ = new_G1766_ & new_G1762_ & new_G1751_;
  assign new_G1785_ = new_G1766_ & new_G1757_ & new_G1754_;
  assign new_G2819_ = ~new_G2817_ | ~new_G2818_;
  assign new_G2824_ = ~new_G2822_ | ~new_G2823_;
  assign new_G4059_ = ~new_G4057_ | ~new_G4058_;
  assign new_G4064_ = ~new_G4062_ | ~new_G4063_;
  assign new_G5081_ = ~new_G5079_ | ~new_G5080_;
  assign new_G5091_ = ~new_G5089_ | ~new_G5090_;
  assign new_G5651_ = ~new_G5649_ | ~new_G5650_;
  assign new_G5661_ = ~new_G5659_ | ~new_G5660_;
  assign new_G6233_ = ~new_G6231_ | ~new_G6232_;
  assign new_G6327_ = ~new_G6321_;
  assign new_G6252_ = ~new_G6321_ | ~new_G6328_;
  assign new_G7107_ = ~new_G7101_;
  assign new_G7110_ = ~new_G7101_ | ~new_G7108_;
  assign new_G7195_ = ~new_G7189_;
  assign new_G7120_ = ~new_G7189_ | ~new_G7196_;
  assign new_G5737_ = new_G1785_ | new_G1784_ | new_G1782_ | new_G1783_;
  assign new_G6251_ = ~new_G6324_ | ~new_G6327_;
  assign new_G7109_ = ~new_G7104_ | ~new_G7107_;
  assign new_G7119_ = ~new_G7192_ | ~new_G7195_;
  assign new_G5087_ = ~new_G5081_;
  assign new_G985_ = ~new_G5081_ | ~new_G5088_;
  assign new_G5097_ = ~new_G5091_;
  assign new_G988_ = ~new_G5091_ | ~new_G5098_;
  assign new_G5657_ = ~new_G5651_;
  assign new_G1776_ = ~new_G5651_ | ~new_G5658_;
  assign new_G5667_ = ~new_G5661_;
  assign new_G1779_ = ~new_G5661_ | ~new_G5668_;
  assign new_G2844_ = new_G2833_ & new_G2824_ & new_G2784_;
  assign new_G2845_ = new_G2833_ & new_G2819_ & new_G2780_;
  assign new_G2846_ = new_G2828_ & new_G2824_ & new_G2813_;
  assign new_G2847_ = new_G2828_ & new_G2819_ & new_G2816_;
  assign new_G4083_ = new_G4072_ & new_G4064_ & new_G4032_;
  assign new_G4084_ = new_G4072_ & new_G4059_ & new_G4028_;
  assign new_G4085_ = new_G4067_ & new_G4064_ & new_G4053_;
  assign new_G4086_ = new_G4067_ & new_G4059_ & new_G4056_;
  assign new_G6239_ = ~new_G6233_;
  assign new_G6242_ = ~new_G6233_ | ~new_G6240_;
  assign new_G6253_ = ~new_G6251_ | ~new_G6252_;
  assign new_G7111_ = ~new_G7109_ | ~new_G7110_;
  assign new_G7121_ = ~new_G7119_ | ~new_G7120_;
  assign new_G984_ = ~new_G5084_ | ~new_G5087_;
  assign new_G987_ = ~new_G5094_ | ~new_G5097_;
  assign new_G1775_ = ~new_G5654_ | ~new_G5657_;
  assign new_G1778_ = ~new_G5664_ | ~new_G5667_;
  assign new_G5743_ = ~new_G5737_;
  assign new_G6241_ = ~new_G6236_ | ~new_G6239_;
  assign new_G6329_ = new_G2847_ | new_G2846_ | new_G2844_ | new_G2845_;
  assign new_G7197_ = new_G4086_ | new_G4085_ | new_G4083_ | new_G4084_;
  assign new_G986_ = ~new_G984_ | ~new_G985_;
  assign new_G989_ = ~new_G987_ | ~new_G988_;
  assign new_G1777_ = ~new_G1775_ | ~new_G1776_;
  assign new_G1780_ = ~new_G1778_ | ~new_G1779_;
  assign new_G6259_ = ~new_G6253_;
  assign new_G2841_ = ~new_G6253_ | ~new_G6260_;
  assign new_G7117_ = ~new_G7111_;
  assign new_G4077_ = ~new_G7111_ | ~new_G7118_;
  assign new_G7127_ = ~new_G7121_;
  assign new_G4080_ = ~new_G7121_ | ~new_G7128_;
  assign new_G6243_ = ~new_G6241_ | ~new_G6242_;
  assign new_G990_ = ~new_G989_;
  assign new_G996_ = new_G975_ & new_G986_;
  assign new_G1781_ = ~new_G1780_;
  assign new_G1787_ = new_G1766_ & new_G1777_;
  assign new_G2840_ = ~new_G6256_ | ~new_G6259_;
  assign new_G6335_ = ~new_G6329_;
  assign new_G4076_ = ~new_G7114_ | ~new_G7117_;
  assign new_G4079_ = ~new_G7124_ | ~new_G7127_;
  assign new_G7203_ = ~new_G7197_;
  assign new_G995_ = new_G990_ & new_G980_;
  assign new_G1786_ = new_G1781_ & new_G1771_;
  assign new_G6249_ = ~new_G6243_;
  assign new_G2838_ = ~new_G6243_ | ~new_G6250_;
  assign new_G2842_ = ~new_G2840_ | ~new_G2841_;
  assign new_G4078_ = ~new_G4076_ | ~new_G4077_;
  assign new_G4081_ = ~new_G4079_ | ~new_G4080_;
  assign new_G2837_ = ~new_G6246_ | ~new_G6249_;
  assign new_G2843_ = ~new_G2842_;
  assign new_G4082_ = ~new_G4081_;
  assign new_G4088_ = new_G4067_ & new_G4078_;
  assign new_G5170_ = new_G995_ | new_G996_;
  assign new_G5740_ = new_G1786_ | new_G1787_;
  assign new_G2839_ = ~new_G2837_ | ~new_G2838_;
  assign new_G2848_ = new_G2843_ & new_G2833_;
  assign new_G4087_ = new_G4082_ & new_G4072_;
  assign new_G1791_ = ~new_G5740_ | ~new_G5743_;
  assign new_G1003_ = ~new_G5170_ | ~new_G5173_;
  assign new_G5174_ = ~new_G5170_;
  assign new_G5744_ = ~new_G5740_;
  assign new_G2849_ = new_G2828_ & new_G2839_;
  assign new_G7200_ = new_G4087_ | new_G4088_;
  assign new_G1792_ = ~new_G5737_ | ~new_G5744_;
  assign new_G1004_ = ~new_G5167_ | ~new_G5174_;
  assign new_G6332_ = new_G2848_ | new_G2849_;
  assign new_G320_ = ~new_G1791_ | ~new_G1792_;
  assign new_G337_ = ~new_G1003_ | ~new_G1004_;
  assign new_G4092_ = ~new_G7200_ | ~new_G7203_;
  assign new_G7204_ = ~new_G7200_;
  assign G321 = ~new_G320_;
  assign G338 = ~new_G337_;
  assign new_G4093_ = ~new_G7197_ | ~new_G7204_;
  assign new_G2855_ = ~new_G6332_ | ~new_G6335_;
  assign new_G6336_ = ~new_G6332_;
  assign new_G369_ = ~new_G4092_ | ~new_G4093_;
  assign new_G2856_ = ~new_G6329_ | ~new_G6336_;
  assign G370 = ~new_G369_;
  assign new_G398_ = ~new_G2855_ | ~new_G2856_;
  assign G399 = ~new_G398_;
endmodule


