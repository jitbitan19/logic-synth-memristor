// NOR_NOT mapped module b10_C

module b10_C (
  input  G_BUTTON,
  input  KEY     ,
  input  START   ,
  input  TEST    ,
  input  RTS     ,
  input  RTR     ,
  input  VOTO0_REG_SCAN_IN,
  input  V_IN_3_ ,
  input  V_IN_2_ ,
  input  V_IN_1_ ,
  input  V_IN_0_ ,
  input  STATO_REG_3__SCAN_IN,
  input  STATO_REG_2__SCAN_IN,
  input  STATO_REG_1__SCAN_IN,
  input  STATO_REG_0__SCAN_IN,
  input  V_OUT_REG_3__SCAN_IN,
  input  V_OUT_REG_2__SCAN_IN,
  input  V_OUT_REG_1__SCAN_IN,
  input  V_OUT_REG_0__SCAN_IN,
  input  SIGN_REG_3__SCAN_IN,
  input  VOTO1_REG_SCAN_IN,
  input  CTR_REG_SCAN_IN,
  input  VOTO3_REG_SCAN_IN,
  input  LAST_R_REG_SCAN_IN,
  input  CTS_REG_SCAN_IN,
  input  VOTO2_REG_SCAN_IN,
  input  LAST_G_REG_SCAN_IN,
  output CTS     ,
  output CTR     ,
  output V_OUT_3_,
  output V_OUT_2_,
  output V_OUT_1_,
  output V_OUT_0_,
  output STATO_REG_3__SCAN_OUT,
  output STATO_REG_2__SCAN_OUT,
  output STATO_REG_1__SCAN_OUT,
  output STATO_REG_0__SCAN_OUT,
  output V_OUT_REG_3__SCAN_OUT,
  output V_OUT_REG_2__SCAN_OUT,
  output V_OUT_REG_1__SCAN_OUT,
  output V_OUT_REG_0__SCAN_OUT,
  output SIGN_REG_3__SCAN_OUT,
  output VOTO1_REG_SCAN_OUT,
  output CTR_REG_SCAN_OUT,
  output VOTO3_REG_SCAN_OUT,
  output LAST_R_REG_SCAN_OUT,
  output CTS_REG_SCAN_OUT,
  output VOTO2_REG_SCAN_OUT,
  output LAST_G_REG_SCAN_OUT,
  output VOTO0_REG_SCAN_OUT);

  wire wr_24;
  wire wr_25;
  wire wr_26;
  wire wr_27;
  wire wr_28;
  wire wr_29;
  wire wr_30;
  wire wr_31;
  wire wr_32;
  wire wr_33;
  wire wr_34;
  wire wr_35;
  wire wr_36;
  wire wr_37;
  wire wr_38;
  wire wr_39;
  wire wr_40;
  wire wr_41;
  wire wr_42;
  wire wr_43;
  wire wr_44;
  wire wr_45;
  wire wr_46;
  wire wr_47;
  wire wr_48;
  wire wr_49;
  wire wr_50;
  wire wr_51;
  wire wr_52;
  wire wr_53;
  wire wr_54;
  wire wr_55;
  wire wr_56;
  wire wr_57;
  wire wr_58;
  wire wr_59;
  wire wr_60;
  wire wr_61;
  wire wr_62;
  wire wr_63;
  wire wr_64;
  wire wr_65;
  wire wr_66;
  wire wr_67;
  wire wr_68;
  wire wr_69;
  wire wr_70;
  wire wr_71;
  wire wr_72;
  wire wr_73;
  wire wr_74;
  wire wr_75;
  wire wr_76;
  wire wr_77;
  wire wr_78;
  wire wr_79;
  wire wr_80;
  wire wr_81;
  wire wr_82;
  wire wr_83;
  wire wr_84;
  wire wr_85;
  wire wr_86;
  wire wr_87;
  wire wr_88;
  wire wr_89;
  wire wr_90;
  wire wr_91;
  wire wr_92;
  wire wr_93;
  wire wr_94;
  wire wr_95;
  wire wr_96;
  wire wr_97;
  wire wr_98;
  wire wr_99;
  wire wr_100;
  wire wr_101;
  wire wr_102;
  wire wr_103;
  wire wr_104;
  wire wr_105;
  wire wr_106;
  wire wr_107;
  wire wr_108;
  wire wr_109;
  wire wr_110;
  wire wr_111;
  wire wr_112;
  wire wr_113;
  wire wr_114;
  wire wr_115;
  wire wr_116;
  wire wr_117;
  wire wr_118;
  wire wr_119;
  wire wr_120;
  wire wr_121;
  wire wr_122;
  wire wr_123;
  wire wr_124;
  wire wr_125;
  wire wr_126;
  wire wr_127;
  wire wr_128;
  wire wr_129;
  wire wr_130;
  wire wr_131;
  wire wr_132;
  wire wr_133;
  wire wr_134;
  wire wr_135;
  wire wr_136;
  wire wr_137;
  wire wr_138;
  wire wr_139;
  wire wr_140;
  wire wr_141;
  wire wr_142;
  wire wr_143;
  wire wr_144;
  wire wr_145;
  wire wr_146;
  wire wr_147;
  wire wr_148;
  wire wr_149;
  wire wr_150;
  wire wr_151;
  wire wr_152;
  wire wr_153;
  wire wr_154;
  wire wr_155;
  wire wr_156;
  wire wr_157;
  wire wr_158;
  wire wr_159;
  wire wr_160;
  wire wr_161;
  wire wr_162;
  wire wr_163;
  wire wr_164;
  wire wr_165;
  wire wr_166;
  wire wr_167;
  wire wr_168;
  wire wr_169;
  wire wr_170;
  wire wr_171;
  wire wr_172;
  wire wr_173;
  wire wr_174;
  wire wr_175;
  wire wr_176;
  wire wr_177;
  wire wr_178;
  wire wr_179;
  wire wr_180;
  wire wr_181;
  wire wr_182;
  wire wr_183;
  wire wr_184;
  wire wr_185;
  wire wr_186;
  wire wr_187;
  wire wr_188;
  wire wr_189;
  wire wr_190;
  wire wr_191;
  wire wr_192;
  wire wr_193;
  wire wr_194;
  wire wr_195;
  wire wr_196;
  wire wr_197;
  wire wr_198;
  wire wr_199;
  wire wr_200;
  wire wr_201;
  wire wr_202;
  wire wr_203;
  wire wr_204;
  wire wr_205;
  wire wr_206;
  wire wr_207;
  wire wr_208;
  wire wr_209;
  wire wr_210;
  wire wr_211;
  wire wr_212;
  wire wr_213;
  wire wr_214;
  wire wr_215;
  wire wr_216;
  wire wr_217;
  wire wr_218;
  wire wr_219;
  wire wr_220;
  wire wr_221;
  wire wr_222;
  wire wr_223;
  wire wr_224;
  wire wr_225;
  wire wr_226;
  wire wr_227;
  wire wr_228;
  wire wr_229;
  wire wr_230;
  wire wr_231;
  wire wr_232;
  wire wr_233;
  wire wr_234;
  wire wr_235;
  wire wr_236;
  wire wr_237;
  wire wr_238;
  wire wr_239;
  wire wr_240;
  wire wr_241;
  wire wr_242;
  wire wr_243;
  wire wr_244;
  wire wr_245;
  wire wr_246;
  wire wr_247;
  wire wr_248;
  wire wr_249;
  wire wr_250;
  wire wr_251;
  wire wr_252;
  wire wr_253;
  wire wr_254;
  wire wr_255;
  wire wr_256;
  wire wr_257;
  wire wr_258;
  wire wr_259;
  wire wr_260;
  wire wr_261;
  wire wr_262;
  wire wr_263;
  wire wr_264;
  wire wr_265;
  wire wr_266;
  wire wr_267;
  wire wr_268;
  wire wr_269;
  wire wr_270;
  wire wr_271;
  wire wr_272;
  wire wr_273;
  wire wr_274;
  wire wr_275;
  wire wr_276;
  wire wr_277;
  wire wr_278;
  wire wr_279;
  wire wr_280;
  wire wr_281;
  wire wr_282;
  wire wr_283;

  not    g1( wr_66   ,           V_IN_3_ );
  not    g2( wr_67   ,           V_IN_2_ );
  nor    g3( wr_75   , STATO_REG_1__SCAN_IN, RTR     );
  not    g4( wr_31   ,           STATO_REG_1__SCAN_IN);
  not    g5( wr_32   ,           STATO_REG_2__SCAN_IN);
  not    g6( wr_45   ,           STATO_REG_0__SCAN_IN);
  not    g7( wr_65   ,           V_IN_0_ );
  nor    g8( wr_25   , STATO_REG_2__SCAN_IN, STATO_REG_3__SCAN_IN);
  not    g9( wr_24   ,           STATO_REG_3__SCAN_IN);
  not   g10( wr_46   ,           START   );
  not   g11( wr_64   ,           V_IN_1_ );
  not   g12( wr_82   ,           RTR     );
  nor   g13( wr_98   , VOTO3_REG_SCAN_IN, VOTO0_REG_SCAN_IN);
  not   g14( wr_30   ,           RTS     );
  not   g15( wr_97   ,           VOTO1_REG_SCAN_IN);
  not   g16( wr_96   ,           VOTO2_REG_SCAN_IN);
  not   g17( wr_157  ,           VOTO0_REG_SCAN_IN);
  not   g18( wr_190  ,           G_BUTTON);
  not   g19( wr_174  ,           KEY     );
  nor   g20( wr_237  , STATO_REG_0__SCAN_IN, STATO_REG_3__SCAN_IN);
  not   g21( wr_143  ,           VOTO3_REG_SCAN_IN);
  not   g22( wr_146  ,           V_OUT_REG_3__SCAN_IN);
  not   g23( wr_150  ,           V_OUT_REG_2__SCAN_IN);
  not   g24( wr_154  ,           V_OUT_REG_1__SCAN_IN);
  not   g25( wr_159  ,           V_OUT_REG_0__SCAN_IN);
  not   g26( wr_163  ,           SIGN_REG_3__SCAN_IN);
  not   g27( wr_201  ,           CTR_REG_SCAN_IN);
  not   g28( wr_236  ,           CTS_REG_SCAN_IN);
  not   g29( wr_267  ,           LAST_G_REG_SCAN_IN);
  not   g30( wr_232  ,           LAST_R_REG_SCAN_IN);
  not   g31( CTS     ,           CTS_REG_SCAN_IN);
  not   g32( CTR     ,           CTR_REG_SCAN_IN);
  not   g33( V_OUT_3_,           V_OUT_REG_3__SCAN_IN);
  not   g34( V_OUT_2_,           V_OUT_REG_2__SCAN_IN);
  not   g35( V_OUT_1_,           V_OUT_REG_1__SCAN_IN);
  not   g36( V_OUT_0_,           V_OUT_REG_0__SCAN_IN);
  nor   g37( wr_68   , wr_67   , wr_66   );
  nor   g38( wr_76   , wr_75   , STATO_REG_0__SCAN_IN);
  nor   g39( wr_33   , STATO_REG_0__SCAN_IN, wr_32   );
  nor   g40( wr_50   , wr_45   , wr_31   );
  nor   g41( wr_74   , wr_31   , STATO_REG_2__SCAN_IN);
  not   g42( wr_26   ,           wr_25   );
  nor   g43( wr_40   , wr_31   , STATO_REG_3__SCAN_IN);
  nor   g44( wr_59   , wr_45   , STATO_REG_1__SCAN_IN);
  nor   g45( wr_61   , wr_32   , RTS     );
  not   g46( wr_99   ,           wr_98   );
  nor   g47( wr_168  , STATO_REG_2__SCAN_IN, wr_24   );
  nor   g48( wr_202  , STATO_REG_1__SCAN_IN, wr_32   );
  nor   g49( wr_115  , wr_45   , STATO_REG_3__SCAN_IN);
  nor   g50( wr_116  , STATO_REG_0__SCAN_IN, wr_24   );
  nor   g51( wr_215  , VOTO2_REG_SCAN_IN, wr_157  );
  nor   g52( wr_216  , wr_96   , VOTO0_REG_SCAN_IN);
  nor   g53( wr_205  , wr_31   , RTS     );
  nor   g54( wr_206  , STATO_REG_1__SCAN_IN, wr_24   );
  nor   g55( wr_240  , STATO_REG_0__SCAN_IN, wr_31   );
  nor   g56( wr_224  , wr_46   , KEY     );
  nor   g57( wr_233  , wr_31   , wr_174  );
  nor   g58( wr_271  , SIGN_REG_3__SCAN_IN, wr_24   );
  nor   g59( wr_238  , wr_237  , wr_82   );
  nor   g60( wr_162  , wr_45   , wr_24   );
  not   g61( wr_69   ,           wr_68   );
  not   g62( wr_77   ,           wr_76   );
  not   g63( wr_34   ,           wr_33   );
  not   g64( wr_51   ,           wr_50   );
  nor   g65( wr_47   , wr_26   , wr_46   );
  not   g66( wr_41   ,           wr_40   );
  nor   g67( wr_27   , wr_26   , STATO_REG_0__SCAN_IN);
  not   g68( wr_60   ,           wr_59   );
  not   g69( wr_62   ,           wr_61   );
  nor   g70( wr_100  , wr_99   , wr_97   );
  not   g71( wr_169  ,           wr_168  );
  nor   g72( wr_203  , wr_202  , wr_74   );
  nor   g73( wr_117  , wr_116  , wr_115  );
  not   g74( wr_175  ,           wr_74   );
  nor   g75( wr_217  , wr_216  , wr_215  );
  nor   g76( wr_207  , wr_206  , wr_205  );
  not   g77( wr_250  ,           wr_206  );
  nor   g78( wr_225  , wr_224  , wr_50   );
  not   g79( wr_234  ,           wr_233  );
  nor   g80( wr_70   , wr_69   , wr_65   );
  nor   g81( wr_78   , wr_77   , wr_74   );
  nor   g82( wr_52   , wr_51   , wr_32   );
  nor   g83( wr_83   , wr_34   , wr_82   );
  not   g84( wr_48   ,           wr_47   );
  nor   g85( wr_35   , wr_34   , wr_31   );
  nor   g86( wr_42   , wr_41   , STATO_REG_2__SCAN_IN);
  not   g87( wr_28   ,           wr_27   );
  nor   g88( wr_63   , wr_62   , wr_60   );
  not   g89( wr_101  ,           wr_100  );
  nor   g90( wr_170  , wr_169  , wr_60   );
  nor   g91( wr_185  , wr_60   , wr_46   );
  not   g92( wr_204  ,           wr_203  );
  not   g93( wr_219  ,           wr_217  );
  nor   g94( wr_276  , wr_117  , wr_175  );
  nor   g95( wr_176  , wr_175  , wr_174  );
  not   g96( wr_208  ,           wr_207  );
  nor   g97( wr_218  , wr_217  , VOTO1_REG_SCAN_IN);
  nor   g98( wr_239  , wr_60   , wr_24   );
  nor   g99( wr_247  , wr_60   , wr_82   );
  nor  g100( wr_251  , wr_250  , wr_34   );
  nor  g101( wr_226  , wr_225  , wr_26   );
  nor  g102( wr_118  , wr_117  , wr_31   );
  nor  g103( wr_125  , wr_41   , STATO_REG_0__SCAN_IN);
  not  g104( wr_71   ,           wr_70   );
  nor  g105( wr_79   , wr_78   , wr_24   );
  not  g106( wr_53   ,           wr_52   );
  not  g107( wr_84   ,           wr_83   );
  nor  g108( wr_49   , wr_48   , wr_45   );
  not  g109( wr_36   ,           wr_35   );
  not  g110( wr_43   ,           wr_42   );
  nor  g111( wr_29   , wr_28   , STATO_REG_1__SCAN_IN);
  nor  g112( wr_102  , wr_101  , wr_96   );
  nor  g113( wr_180  , wr_28   , wr_46   );
  not  g114( wr_186  ,           wr_185  );
  nor  g115( wr_241  , wr_240  , wr_204  );
  nor  g116( wr_95   , wr_28   , TEST    );
  nor  g117( wr_220  , wr_219  , wr_97   );
  nor  g118( wr_272  , wr_28   , wr_174  );
  not  g119( wr_177  ,           wr_176  );
  nor  g120( wr_209  , wr_208  , STATO_REG_0__SCAN_IN);
  not  g121( wr_248  ,           wr_247  );
  nor  g122( wr_72   , wr_71   , wr_64   );
  not  g123( wr_80   ,           wr_79   );
  nor  g124( wr_54   , wr_53   , RTR     );
  nor  g125( wr_85   , wr_84   , STATO_REG_1__SCAN_IN);
  nor  g126( wr_37   , wr_36   , wr_30   );
  nor  g127( wr_44   , wr_43   , START   );
  not  g128( wr_103  ,           wr_102  );
  not  g129( wr_181  ,           wr_180  );
  nor  g130( wr_187  , wr_186  , STATO_REG_2__SCAN_IN);
  nor  g131( wr_110  , wr_102  , STATO_REG_0__SCAN_IN);
  nor  g132( wr_171  , wr_36   , STATO_REG_3__SCAN_IN);
  not  g133( wr_242  ,           wr_241  );
  nor  g134( wr_221  , wr_220  , wr_218  );
  nor  g135( wr_273  , wr_272  , wr_271  );
  not  g136( wr_164  ,           wr_95   );
  nor  g137( wr_178  , wr_177  , VOTO1_REG_SCAN_IN);
  not  g138( wr_210  ,           wr_209  );
  nor  g139( wr_249  , wr_248  , wr_26   );
  nor  g140( wr_258  , wr_177  , VOTO2_REG_SCAN_IN);
  nor  g141( wr_73   , wr_72   , wr_45   );
  nor  g142( wr_55   , wr_54   , wr_49   );
  nor  g143( wr_38   , wr_37   , wr_29   );
  nor  g144( wr_133  , wr_103  , STATO_REG_3__SCAN_IN);
  nor  g145( wr_191  , wr_181  , wr_190  );
  nor  g146( wr_104  , wr_103  , wr_34   );
  nor  g147( wr_172  , wr_171  , wr_170  );
  nor  g148( wr_182  , wr_181  , KEY     );
  nor  g149( wr_243  , wr_242  , wr_239  );
  nor  g150( wr_252  , wr_251  , wr_85   );
  nor  g151( wr_222  , wr_221  , wr_51   );
  nor  g152( wr_235  , wr_234  , wr_181  );
  nor  g153( wr_274  , wr_273  , wr_31   );
  not  g154( wr_144  ,           wr_85   );
  nor  g155( wr_165  , wr_164  , STATO_REG_1__SCAN_IN);
  nor  g156( wr_211  , wr_210  , wr_204  );
  nor  g157( wr_147  , wr_85   , wr_146  );
  nor  g158( wr_151  , wr_85   , wr_150  );
  nor  g159( wr_155  , wr_85   , wr_154  );
  nor  g160( wr_160  , wr_85   , wr_159  );
  nor  g161( wr_81   , wr_80   , wr_73   );
  not  g162( wr_56   ,           wr_55   );
  not  g163( wr_39   ,           wr_38   );
  nor  g164( wr_134  , wr_133  , STATO_REG_0__SCAN_IN);
  not  g165( wr_192  ,           wr_191  );
  nor  g166( wr_105  , wr_104  , wr_95   );
  nor  g167( wr_173  , wr_172  , wr_64   );
  nor  g168( wr_214  , wr_172  , wr_66   );
  not  g169( wr_244  ,           wr_243  );
  not  g170( wr_253  ,           wr_252  );
  nor  g171( wr_257  , wr_172  , wr_67   );
  nor  g172( wr_270  , wr_172  , wr_65   );
  not  g173( wr_265  ,           wr_235  );
  nor  g174( wr_145  , wr_144  , wr_143  );
  nor  g175( wr_149  , wr_144  , wr_96   );
  nor  g176( wr_153  , wr_144  , wr_97   );
  nor  g177( wr_158  , wr_144  , wr_157  );
  nor  g178( wr_166  , wr_165  , wr_163  );
  nor  g179( wr_212  , wr_211  , wr_201  );
  nor  g180( wr_268  , wr_235  , wr_267  );
  nor  g181( LAST_R_REG_SCAN_OUT, wr_235  , wr_232  );
  nor  g182( wr_86   , wr_85   , wr_81   );
  nor  g183( wr_57   , wr_56   , wr_44   );
  nor  g184( wr_183  , wr_170  , wr_39   );
  not  g185( wr_135  ,           wr_134  );
  nor  g186( wr_193  , wr_192  , LAST_G_REG_SCAN_IN);
  nor  g187( wr_179  , wr_178  , wr_173  );
  nor  g188( wr_223  , wr_222  , wr_214  );
  nor  g189( wr_245  , wr_244  , wr_238  );
  nor  g190( wr_254  , wr_253  , wr_249  );
  nor  g191( wr_259  , wr_258  , wr_257  );
  nor  g192( wr_275  , wr_274  , wr_270  );
  nor  g193( wr_266  , wr_265  , wr_190  );
  nor  g194( wr_148  , wr_147  , wr_145  );
  nor  g195( wr_152  , wr_151  , wr_149  );
  nor  g196( wr_156  , wr_155  , wr_153  );
  nor  g197( wr_161  , wr_160  , wr_158  );
  nor  g198( wr_167  , wr_166  , wr_162  );
  nor  g199( wr_213  , wr_212  , wr_63   );
  not  g200( wr_87   ,           wr_86   );
  not  g201( wr_58   ,           wr_57   );
  not  g202( wr_184  ,           wr_183  );
  nor  g203( wr_136  , wr_135  , STATO_REG_1__SCAN_IN);
  nor  g204( wr_246  , wr_245  , wr_236  );
  not  g205( wr_255  ,           wr_254  );
  nor  g206( wr_269  , wr_268  , wr_266  );
  not  g207( V_OUT_REG_3__SCAN_OUT,           wr_148  );
  not  g208( V_OUT_REG_2__SCAN_OUT,           wr_152  );
  not  g209( V_OUT_REG_1__SCAN_OUT,           wr_156  );
  not  g210( V_OUT_REG_0__SCAN_OUT,           wr_161  );
  not  g211( SIGN_REG_3__SCAN_OUT,           wr_167  );
  not  g212( CTR_REG_SCAN_OUT,           wr_213  );
  nor  g213( wr_88   , wr_87   , wr_63   );
  nor  g214( wr_188  , wr_187  , wr_184  );
  nor  g215( wr_277  , wr_276  , wr_184  );
  nor  g216( wr_137  , wr_136  , wr_35   );
  nor  g217( wr_256  , wr_255  , wr_246  );
  not  g218( LAST_G_REG_SCAN_OUT,           wr_269  );
  not  g219( wr_89   ,           wr_88   );
  not  g220( wr_189  ,           wr_188  );
  not  g221( wr_278  ,           wr_277  );
  not  g222( wr_138  ,           wr_137  );
  not  g223( CTS_REG_SCAN_OUT,           wr_256  );
  nor  g224( wr_90   , wr_89   , wr_58   );
  nor  g225( wr_194  , wr_193  , wr_189  );
  nor  g226( wr_227  , wr_226  , wr_189  );
  nor  g227( wr_260  , wr_189  , wr_182  );
  nor  g228( wr_279  , wr_278  , wr_47   );
  nor  g229( wr_139  , wr_138  , wr_27   );
  not  g230( wr_91   ,           wr_90   );
  not  g231( wr_195  ,           wr_194  );
  not  g232( wr_229  ,           wr_227  );
  not  g233( wr_262  ,           wr_260  );
  not  g234( wr_281  ,           wr_279  );
  nor  g235( wr_228  , wr_227  , wr_223  );
  nor  g236( wr_261  , wr_260  , wr_259  );
  nor  g237( wr_280  , wr_279  , wr_275  );
  nor  g238( wr_92   , wr_91   , wr_39   );
  nor  g239( wr_196  , wr_195  , wr_182  );
  nor  g240( wr_230  , wr_229  , wr_143  );
  nor  g241( wr_263  , wr_262  , wr_96   );
  nor  g242( wr_282  , wr_281  , wr_157  );
  nor  g243( wr_111  , wr_110  , wr_92   );
  not  g244( wr_126  ,           wr_92   );
  nor  g245( wr_106  , wr_105  , wr_92   );
  nor  g246( wr_122  , wr_92   , wr_45   );
  nor  g247( wr_93   , wr_92   , STATO_REG_0__SCAN_IN);
  not  g248( wr_198  ,           wr_196  );
  nor  g249( wr_140  , wr_139  , wr_92   );
  nor  g250( wr_197  , wr_196  , wr_179  );
  nor  g251( wr_231  , wr_230  , wr_228  );
  nor  g252( wr_264  , wr_263  , wr_261  );
  nor  g253( wr_283  , wr_282  , wr_280  );
  not  g254( wr_112  ,           wr_111  );
  nor  g255( wr_127  , wr_126  , wr_31   );
  not  g256( wr_107  ,           wr_106  );
  not  g257( wr_123  ,           wr_122  );
  nor  g258( wr_94   , wr_93   , wr_24   );
  nor  g259( wr_141  , wr_126  , wr_45   );
  nor  g260( wr_199  , wr_198  , wr_97   );
  not  g261( VOTO3_REG_SCAN_OUT,           wr_231  );
  not  g262( VOTO2_REG_SCAN_OUT,           wr_264  );
  not  g263( VOTO0_REG_SCAN_OUT,           wr_283  );
  nor  g264( wr_113  , wr_112  , wr_59   );
  nor  g265( wr_128  , wr_127  , wr_35   );
  nor  g266( wr_108  , wr_107  , STATO_REG_1__SCAN_IN);
  nor  g267( wr_124  , wr_123  , wr_40   );
  nor  g268( wr_142  , wr_141  , wr_140  );
  nor  g269( wr_200  , wr_199  , wr_197  );
  nor  g270( wr_114  , wr_113  , wr_32   );
  not  g271( wr_129  ,           wr_128  );
  nor  g272( wr_109  , wr_108  , wr_94   );
  not  g273( STATO_REG_0__SCAN_OUT,           wr_142  );
  not  g274( VOTO1_REG_SCAN_OUT,           wr_200  );
  nor  g275( wr_119  , wr_118  , wr_114  );
  nor  g276( wr_130  , wr_129  , wr_125  );
  not  g277( STATO_REG_3__SCAN_OUT,           wr_109  );
  not  g278( wr_120  ,           wr_119  );
  not  g279( wr_131  ,           wr_130  );
  nor  g280( wr_121  , wr_120  , wr_35   );
  nor  g281( wr_132  , wr_131  , wr_124  );
  not  g282( STATO_REG_2__SCAN_OUT,           wr_121  );
  not  g283( STATO_REG_1__SCAN_OUT,           wr_132  );

endmodule
