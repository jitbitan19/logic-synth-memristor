// NOR_NOT mapped module c880

module c880 (
  input  G1gat   ,
  input  G8gat   ,
  input  G13gat  ,
  input  G17gat  ,
  input  G26gat  ,
  input  G29gat  ,
  input  G36gat  ,
  input  G42gat  ,
  input  G51gat  ,
  input  G55gat  ,
  input  G59gat  ,
  input  G68gat  ,
  input  G72gat  ,
  input  G73gat  ,
  input  G74gat  ,
  input  G75gat  ,
  input  G80gat  ,
  input  G85gat  ,
  input  G86gat  ,
  input  G87gat  ,
  input  G88gat  ,
  input  G89gat  ,
  input  G90gat  ,
  input  G91gat  ,
  input  G96gat  ,
  input  G101gat ,
  input  G106gat ,
  input  G111gat ,
  input  G116gat ,
  input  G121gat ,
  input  G126gat ,
  input  G130gat ,
  input  G135gat ,
  input  G138gat ,
  input  G143gat ,
  input  G146gat ,
  input  G149gat ,
  input  G152gat ,
  input  G153gat ,
  input  G156gat ,
  input  G159gat ,
  input  G165gat ,
  input  G171gat ,
  input  G177gat ,
  input  G183gat ,
  input  G189gat ,
  input  G195gat ,
  input  G201gat ,
  input  G207gat ,
  input  G210gat ,
  input  G219gat ,
  input  G228gat ,
  input  G237gat ,
  input  G246gat ,
  input  G255gat ,
  input  G259gat ,
  input  G260gat ,
  input  G261gat ,
  input  G267gat ,
  input  G268gat ,
  output G388gat ,
  output G389gat ,
  output G390gat ,
  output G391gat ,
  output G418gat ,
  output G419gat ,
  output G420gat ,
  output G421gat ,
  output G422gat ,
  output G423gat ,
  output G446gat ,
  output G447gat ,
  output G448gat ,
  output G449gat ,
  output G450gat ,
  output G767gat ,
  output G768gat ,
  output G850gat ,
  output G863gat ,
  output G864gat ,
  output G865gat ,
  output G866gat ,
  output G874gat ,
  output G878gat ,
  output G879gat ,
  output G880gat );

  wire wr_27;
  wire wr_28;
  wire wr_29;
  wire wr_30;
  wire wr_31;
  wire wr_32;
  wire wr_33;
  wire wr_34;
  wire wr_35;
  wire wr_36;
  wire wr_37;
  wire wr_38;
  wire wr_39;
  wire wr_40;
  wire wr_41;
  wire wr_42;
  wire wr_43;
  wire wr_44;
  wire wr_45;
  wire wr_46;
  wire wr_47;
  wire wr_48;
  wire wr_49;
  wire wr_50;
  wire wr_51;
  wire wr_52;
  wire wr_53;
  wire wr_54;
  wire wr_55;
  wire wr_56;
  wire wr_57;
  wire wr_58;
  wire wr_59;
  wire wr_60;
  wire wr_61;
  wire wr_62;
  wire wr_63;
  wire wr_64;
  wire wr_65;
  wire wr_66;
  wire wr_67;
  wire wr_68;
  wire wr_69;
  wire wr_70;
  wire wr_71;
  wire wr_72;
  wire wr_73;
  wire wr_74;
  wire wr_75;
  wire wr_76;
  wire wr_77;
  wire wr_78;
  wire wr_79;
  wire wr_80;
  wire wr_81;
  wire wr_82;
  wire wr_83;
  wire wr_84;
  wire wr_85;
  wire wr_86;
  wire wr_87;
  wire wr_88;
  wire wr_89;
  wire wr_90;
  wire wr_91;
  wire wr_92;
  wire wr_93;
  wire wr_94;
  wire wr_95;
  wire wr_96;
  wire wr_97;
  wire wr_98;
  wire wr_99;
  wire wr_100;
  wire wr_101;
  wire wr_102;
  wire wr_103;
  wire wr_104;
  wire wr_105;
  wire wr_106;
  wire wr_107;
  wire wr_108;
  wire wr_109;
  wire wr_110;
  wire wr_111;
  wire wr_112;
  wire wr_113;
  wire wr_114;
  wire wr_115;
  wire wr_116;
  wire wr_117;
  wire wr_118;
  wire wr_119;
  wire wr_120;
  wire wr_121;
  wire wr_122;
  wire wr_123;
  wire wr_124;
  wire wr_125;
  wire wr_126;
  wire wr_127;
  wire wr_128;
  wire wr_129;
  wire wr_130;
  wire wr_131;
  wire wr_132;
  wire wr_133;
  wire wr_134;
  wire wr_135;
  wire wr_136;
  wire wr_137;
  wire wr_138;
  wire wr_139;
  wire wr_140;
  wire wr_141;
  wire wr_142;
  wire wr_143;
  wire wr_144;
  wire wr_145;
  wire wr_146;
  wire wr_147;
  wire wr_148;
  wire wr_149;
  wire wr_150;
  wire wr_151;
  wire wr_152;
  wire wr_153;
  wire wr_154;
  wire wr_155;
  wire wr_156;
  wire wr_157;
  wire wr_158;
  wire wr_159;
  wire wr_160;
  wire wr_161;
  wire wr_162;
  wire wr_163;
  wire wr_164;
  wire wr_165;
  wire wr_166;
  wire wr_167;
  wire wr_168;
  wire wr_169;
  wire wr_170;
  wire wr_171;
  wire wr_172;
  wire wr_173;
  wire wr_174;
  wire wr_175;
  wire wr_176;
  wire wr_177;
  wire wr_178;
  wire wr_179;
  wire wr_180;
  wire wr_181;
  wire wr_182;
  wire wr_183;
  wire wr_184;
  wire wr_185;
  wire wr_186;
  wire wr_187;
  wire wr_188;
  wire wr_189;
  wire wr_190;
  wire wr_191;
  wire wr_192;
  wire wr_193;
  wire wr_194;
  wire wr_195;
  wire wr_196;
  wire wr_197;
  wire wr_198;
  wire wr_199;
  wire wr_200;
  wire wr_201;
  wire wr_202;
  wire wr_203;
  wire wr_204;
  wire wr_205;
  wire wr_206;
  wire wr_207;
  wire wr_208;
  wire wr_209;
  wire wr_210;
  wire wr_211;
  wire wr_212;
  wire wr_213;
  wire wr_214;
  wire wr_215;
  wire wr_216;
  wire wr_217;
  wire wr_218;
  wire wr_219;
  wire wr_220;
  wire wr_221;
  wire wr_222;
  wire wr_223;
  wire wr_224;
  wire wr_225;
  wire wr_226;
  wire wr_227;
  wire wr_228;
  wire wr_229;
  wire wr_230;
  wire wr_231;
  wire wr_232;
  wire wr_233;
  wire wr_234;
  wire wr_235;
  wire wr_236;
  wire wr_237;
  wire wr_238;
  wire wr_239;
  wire wr_240;
  wire wr_241;
  wire wr_242;
  wire wr_243;
  wire wr_244;
  wire wr_245;
  wire wr_246;
  wire wr_247;
  wire wr_248;
  wire wr_249;
  wire wr_250;
  wire wr_251;
  wire wr_252;
  wire wr_253;
  wire wr_254;
  wire wr_255;
  wire wr_256;
  wire wr_257;
  wire wr_258;
  wire wr_259;
  wire wr_260;
  wire wr_261;
  wire wr_262;
  wire wr_263;
  wire wr_264;
  wire wr_265;
  wire wr_266;
  wire wr_267;
  wire wr_268;
  wire wr_269;
  wire wr_270;
  wire wr_271;
  wire wr_272;
  wire wr_273;
  wire wr_274;
  wire wr_275;
  wire wr_276;
  wire wr_277;
  wire wr_278;
  wire wr_279;
  wire wr_280;
  wire wr_281;
  wire wr_282;
  wire wr_283;
  wire wr_284;
  wire wr_285;
  wire wr_286;
  wire wr_287;
  wire wr_288;
  wire wr_289;
  wire wr_290;
  wire wr_291;
  wire wr_292;
  wire wr_293;
  wire wr_294;
  wire wr_295;
  wire wr_296;
  wire wr_297;
  wire wr_298;
  wire wr_299;
  wire wr_300;
  wire wr_301;
  wire wr_302;
  wire wr_303;
  wire wr_304;
  wire wr_305;
  wire wr_306;
  wire wr_307;
  wire wr_308;
  wire wr_309;
  wire wr_310;
  wire wr_311;
  wire wr_312;
  wire wr_313;
  wire wr_314;
  wire wr_315;
  wire wr_316;
  wire wr_317;
  wire wr_318;
  wire wr_319;
  wire wr_320;
  wire wr_321;
  wire wr_322;
  wire wr_323;
  wire wr_324;
  wire wr_325;
  wire wr_326;
  wire wr_327;
  wire wr_328;
  wire wr_329;
  wire wr_330;
  wire wr_331;
  wire wr_332;
  wire wr_333;
  wire wr_334;
  wire wr_335;
  wire wr_336;
  wire wr_337;
  wire wr_338;
  wire wr_339;
  wire wr_340;
  wire wr_341;
  wire wr_342;
  wire wr_343;
  wire wr_344;
  wire wr_345;
  wire wr_346;
  wire wr_347;
  wire wr_348;
  wire wr_349;
  wire wr_350;
  wire wr_351;
  wire wr_352;
  wire wr_353;
  wire wr_354;
  wire wr_355;
  wire wr_356;
  wire wr_357;
  wire wr_358;
  wire wr_359;
  wire wr_360;
  wire wr_361;
  wire wr_362;
  wire wr_363;
  wire wr_364;
  wire wr_365;
  wire wr_366;
  wire wr_367;
  wire wr_368;
  wire wr_369;
  wire wr_370;
  wire wr_371;
  wire wr_372;
  wire wr_373;
  wire wr_374;
  wire wr_375;
  wire wr_376;
  wire wr_377;
  wire wr_378;
  wire wr_379;
  wire wr_380;
  wire wr_381;
  wire wr_382;
  wire wr_383;
  wire wr_384;
  wire wr_385;
  wire wr_386;
  wire wr_387;
  wire wr_388;
  wire wr_389;
  wire wr_390;
  wire wr_391;
  wire wr_392;
  wire wr_393;
  wire wr_394;
  wire wr_395;
  wire wr_396;
  wire wr_397;
  wire wr_398;
  wire wr_399;
  wire wr_400;
  wire wr_401;
  wire wr_402;
  wire wr_403;
  wire wr_404;
  wire wr_405;
  wire wr_406;
  wire wr_407;
  wire wr_408;
  wire wr_409;
  wire wr_410;
  wire wr_411;
  wire wr_412;
  wire wr_413;
  wire wr_414;
  wire wr_415;
  wire wr_416;
  wire wr_417;
  wire wr_418;
  wire wr_419;
  wire wr_420;
  wire wr_421;
  wire wr_422;
  wire wr_423;
  wire wr_424;
  wire wr_425;
  wire wr_426;
  wire wr_427;
  wire wr_428;
  wire wr_429;
  wire wr_430;
  wire wr_431;
  wire wr_432;
  wire wr_433;
  wire wr_434;
  wire wr_435;
  wire wr_436;
  wire wr_437;
  wire wr_438;
  wire wr_439;
  wire wr_440;
  wire wr_441;
  wire wr_442;
  wire wr_443;
  wire wr_444;
  wire wr_445;
  wire wr_446;
  wire wr_447;
  wire wr_448;
  wire wr_449;
  wire wr_450;
  wire wr_451;
  wire wr_452;
  wire wr_453;
  wire wr_454;
  wire wr_455;
  wire wr_456;
  wire wr_457;
  wire wr_458;
  wire wr_459;
  wire wr_460;
  wire wr_461;
  wire wr_462;
  wire wr_463;
  wire wr_464;
  wire wr_465;
  wire wr_466;
  wire wr_467;
  wire wr_468;
  wire wr_469;
  wire wr_470;
  wire wr_471;
  wire wr_472;
  wire wr_473;
  wire wr_474;
  wire wr_475;
  wire wr_476;
  wire wr_477;
  wire wr_478;
  wire wr_479;
  wire wr_480;
  wire wr_481;
  wire wr_482;
  wire wr_483;
  wire wr_484;
  wire wr_485;
  wire wr_486;
  wire wr_487;
  wire wr_488;
  wire wr_489;
  wire wr_490;
  wire wr_491;
  wire wr_492;
  wire wr_493;
  wire wr_494;
  wire wr_495;
  wire wr_496;
  wire wr_497;
  wire wr_498;
  wire wr_499;
  wire wr_500;
  wire wr_501;
  wire wr_502;
  wire wr_503;
  wire wr_504;
  wire wr_505;
  wire wr_506;
  wire wr_507;
  wire wr_508;
  wire wr_509;
  wire wr_510;
  wire wr_511;
  wire wr_512;
  wire wr_513;
  wire wr_514;
  wire wr_515;
  wire wr_516;
  wire wr_517;
  wire wr_518;
  wire wr_519;
  wire wr_520;
  wire wr_521;
  wire wr_522;
  wire wr_523;
  wire wr_524;
  wire wr_525;
  wire wr_526;
  wire wr_527;
  wire wr_528;
  wire wr_529;
  wire wr_530;
  wire wr_531;
  wire wr_532;
  wire wr_533;
  wire wr_534;
  wire wr_535;
  wire wr_536;
  wire wr_537;
  wire wr_538;
  wire wr_539;
  wire wr_540;
  wire wr_541;
  wire wr_542;
  wire wr_543;
  wire wr_544;
  wire wr_545;
  wire wr_546;
  wire wr_547;
  wire wr_548;
  wire wr_549;
  wire wr_550;
  wire wr_551;
  wire wr_552;
  wire wr_553;

  not    g1( wr_27   ,           G75gat  );
  not    g2( wr_28   ,           G29gat  );
  not    g3( wr_29   ,           G42gat  );
  not    g4( wr_33   ,           G80gat  );
  not    g5( wr_38   ,           G8gat   );
  not    g6( wr_39   ,           G1gat   );
  not    g7( wr_41   ,           G17gat  );
  not    g8( wr_46   ,           G26gat  );
  not    g9( wr_50   ,           G59gat  );
  not   g10( wr_62   ,           G51gat  );
  not   g11( wr_65   ,           G55gat  );
  not   g12( wr_102  ,           G111gat );
  not   g13( wr_103  ,           G116gat );
  not   g14( wr_108  ,           G126gat );
  not   g15( wr_151  ,           G201gat );
  not   g16( wr_177  ,           G153gat );
  not   g17( wr_178  ,           G156gat );
  nor   g18( wr_185  , G42gat  , G17gat  );
  not   g19( wr_222  ,           G261gat );
  not   g20( wr_254  ,           G143gat );
  not   g21( wr_275  ,           G146gat );
  not   g22( wr_88   ,           G106gat );
  not   g23( wr_107  ,           G121gat );
  not   g24( wr_146  ,           G189gat );
  not   g25( wr_150  ,           G195gat );
  not   g26( wr_283  ,           G149gat );
  not   g27( wr_380  ,           G138gat );
  not   g28( wr_425  ,           G152gat );
  not   g29( wr_83   ,           G96gat  );
  not   g30( wr_87   ,           G101gat );
  not   g31( wr_145  ,           G183gat );
  not   g32( wr_131  ,           G177gat );
  not   g33( wr_82   ,           G91gat  );
  not   g34( wr_40   ,           G13gat  );
  not   g35( wr_72   ,           G68gat  );
  not   g36( wr_230  ,           G72gat  );
  not   g37( wr_126  ,           G165gat );
  not   g38( wr_130  ,           G171gat );
  not   g39( wr_125  ,           G159gat );
  nor   g40( wr_85   , G96gat  , G91gat  );
  nor   g41( wr_90   , G106gat , G101gat );
  nor   g42( wr_105  , G116gat , G111gat );
  nor   g43( wr_110  , G126gat , G121gat );
  nor   g44( wr_128  , G165gat , G159gat );
  nor   g45( wr_133  , G177gat , G171gat );
  nor   g46( wr_148  , G189gat , G183gat );
  nor   g47( wr_153  , G201gat , G195gat );
  not   g48( wr_229  ,           G73gat  );
  not   g49( wr_242  ,           G255gat );
  not   g50( wr_243  ,           G267gat );
  not   g51( wr_245  ,           G246gat );
  not   g52( wr_343  ,           G259gat );
  not   g53( wr_370  ,           G260gat );
  not   g54( wr_218  ,           G210gat );
  not   g55( wr_220  ,           G219gat );
  not   g56( wr_488  ,           G268gat );
  not   g57( wr_75   ,           G74gat  );
  not   g58( wr_81   ,           G130gat );
  not   g59( wr_101  ,           G135gat );
  not   g60( wr_144  ,           G207gat );
  not   g61( wr_168  ,           G228gat );
  not   g62( wr_213  ,           G237gat );
  not   g63( wr_32   ,           G36gat  );
  not   g64( wr_36   ,           G85gat  );
  not   g65( wr_37   ,           G86gat  );
  not   g66( wr_58   ,           G90gat  );
  nor   g67( wr_59   , G88gat  , G87gat  );
  not   g68( wr_80   ,           G89gat  );
  nor   g69( wr_34   , wr_33   , wr_28   );
  nor   g70( wr_55   , wr_50   , wr_29   );
  nor   g71( wr_63   , wr_62   , wr_39   );
  nor   g72( wr_179  , wr_178  , wr_50   );
  nor   g73( wr_186  , wr_29   , wr_41   );
  nor   g74( wr_194  , wr_62   , wr_41   );
  nor   g75( wr_426  , wr_425  , wr_380  );
  nor   g76( wr_399  , wr_380  , wr_62   );
  nor   g77( wr_409  , wr_380  , wr_41   );
  nor   g78( wr_381  , wr_380  , wr_38   );
  nor   g79( wr_66   , wr_65   , wr_40   );
  nor   g80( wr_231  , wr_230  , wr_72   );
  nor   g81( wr_84   , wr_83   , wr_82   );
  nor   g82( wr_89   , wr_88   , wr_87   );
  nor   g83( wr_104  , wr_103  , wr_102  );
  nor   g84( wr_109  , wr_108  , wr_107  );
  nor   g85( wr_127  , wr_126  , wr_125  );
  nor   g86( wr_132  , wr_131  , wr_130  );
  nor   g87( wr_147  , wr_146  , wr_145  );
  nor   g88( wr_152  , wr_151  , wr_150  );
  nor   g89( wr_244  , wr_243  , wr_242  );
  nor   g90( wr_344  , wr_343  , wr_242  );
  nor   g91( wr_371  , wr_370  , wr_242  );
  nor   g92( wr_42   , wr_41   , wr_40   );
  nor   g93( wr_219  , wr_218  , wr_107  );
  nor   g94( wr_274  , wr_218  , wr_88   );
  nor   g95( wr_326  , wr_218  , wr_102  );
  nor   g96( wr_359  , wr_218  , wr_103  );
  nor   g97( wr_465  , wr_218  , wr_87   );
  nor   g98( wr_489  , wr_488  , wr_218  );
  nor   g99( wr_512  , wr_218  , wr_82   );
  nor  g100( wr_541  , wr_218  , wr_83   );
  nor  g101( wr_30   , wr_29   , wr_28   );
  nor  g102( wr_76   , wr_75   , wr_50   );
  nor  g103( wr_51   , wr_33   , wr_50   );
  nor  g104( wr_73   , wr_72   , wr_28   );
  nor  g105( G391gat , wr_37   , wr_36   );
  nor  g106( G423gat , wr_59   , wr_58   );
  nor  g107( G450gat , wr_59   , wr_80   );
  not  g108( wr_35   ,           wr_34   );
  not  g109( wr_56   ,           wr_55   );
  not  g110( wr_64   ,           wr_63   );
  nor  g111( wr_187  , wr_186  , wr_185  );
  not  g112( wr_195  ,           wr_194  );
  nor  g113( wr_385  , wr_179  , wr_65   );
  not  g114( wr_67   ,           wr_66   );
  not  g115( wr_232  ,           wr_231  );
  nor  g116( wr_86   , wr_85   , wr_84   );
  nor  g117( wr_91   , wr_90   , wr_89   );
  nor  g118( wr_106  , wr_105  , wr_104  );
  nor  g119( wr_111  , wr_110  , wr_109  );
  nor  g120( wr_129  , wr_128  , wr_127  );
  nor  g121( wr_134  , wr_133  , wr_132  );
  nor  g122( wr_149  , wr_148  , wr_147  );
  nor  g123( wr_154  , wr_153  , wr_152  );
  not  g124( wr_43   ,           wr_42   );
  not  g125( wr_31   ,           wr_30   );
  not  g126( wr_77   ,           wr_76   );
  not  g127( wr_52   ,           wr_51   );
  not  g128( wr_74   ,           wr_73   );
  nor  g129( G447gat , wr_64   , wr_46   );
  nor  g130( wr_169  , wr_35   , wr_27   );
  not  g131( wr_188  ,           wr_187  );
  nor  g132( wr_196  , wr_195  , wr_39   );
  nor  g133( wr_200  , wr_56   , wr_27   );
  not  g134( wr_386  ,           wr_385  );
  nor  g135( wr_68   , wr_67   , wr_39   );
  nor  g136( wr_233  , wr_232  , wr_50   );
  not  g137( wr_93   ,           wr_86   );
  not  g138( wr_94   ,           wr_91   );
  not  g139( wr_113  ,           wr_106  );
  not  g140( wr_114  ,           wr_111  );
  not  g141( wr_136  ,           wr_129  );
  not  g142( wr_137  ,           wr_134  );
  not  g143( wr_156  ,           wr_149  );
  not  g144( wr_157  ,           wr_154  );
  nor  g145( wr_92   , wr_91   , wr_86   );
  nor  g146( wr_112  , wr_111  , wr_106  );
  nor  g147( wr_135  , wr_134  , wr_129  );
  nor  g148( wr_155  , wr_154  , wr_149  );
  nor  g149( wr_44   , wr_43   , wr_39   );
  nor  g150( G390gat , wr_31   , wr_32   );
  nor  g151( wr_78   , wr_77   , wr_72   );
  nor  g152( wr_53   , wr_52   , wr_27   );
  nor  g153( wr_54   , wr_52   , wr_32   );
  nor  g154( wr_57   , wr_56   , wr_32   );
  nor  g155( G388gat , wr_31   , wr_27   );
  nor  g156( G389gat , wr_35   , wr_32   );
  not  g157( wr_170  ,           wr_169  );
  not  g158( wr_171  ,           G447gat );
  not  g159( wr_197  ,           wr_196  );
  not  g160( wr_69   ,           wr_68   );
  not  g161( wr_234  ,           wr_233  );
  nor  g162( wr_95   , wr_94   , wr_93   );
  nor  g163( wr_115  , wr_114  , wr_113  );
  nor  g164( wr_138  , wr_137  , wr_136  );
  nor  g165( wr_158  , wr_157  , wr_156  );
  not  g166( wr_45   ,           wr_44   );
  not  g167( wr_60   ,           G390gat );
  not  g168( wr_79   ,           wr_78   );
  not  g169( G420gat ,           wr_53   );
  not  g170( G421gat ,           wr_54   );
  not  g171( G422gat ,           wr_57   );
  nor  g172( wr_172  , wr_171  , wr_65   );
  nor  g173( wr_180  , wr_171  , wr_41   );
  nor  g174( wr_189  , wr_171  , wr_178  );
  nor  g175( wr_198  , wr_197  , wr_38   );
  nor  g176( wr_387  , wr_386  , wr_171  );
  nor  g177( wr_390  , wr_170  , wr_171  );
  nor  g178( wr_70   , wr_69   , wr_38   );
  nor  g179( wr_235  , wr_234  , wr_29   );
  nor  g180( wr_96   , wr_95   , wr_92   );
  nor  g181( wr_116  , wr_115  , wr_112  );
  nor  g182( wr_139  , wr_138  , wr_135  );
  nor  g183( wr_159  , wr_158  , wr_155  );
  nor  g184( wr_47   , wr_45   , wr_46   );
  nor  g185( G418gat , wr_45   , wr_38   );
  not  g186( wr_173  ,           wr_172  );
  not  g187( wr_181  ,           wr_180  );
  not  g188( wr_190  ,           wr_189  );
  not  g189( wr_199  ,           wr_198  );
  not  g190( wr_391  ,           wr_390  );
  not  g191( wr_388  ,           wr_387  );
  not  g192( wr_71   ,           wr_70   );
  not  g193( wr_236  ,           wr_235  );
  not  g194( wr_97   ,           wr_96   );
  not  g195( wr_117  ,           wr_116  );
  not  g196( wr_140  ,           wr_139  );
  not  g197( wr_160  ,           wr_159  );
  nor  g198( wr_99   , wr_96   , G130gat );
  nor  g199( wr_119  , wr_116  , G135gat );
  nor  g200( wr_142  , wr_139  , G130gat );
  nor  g201( wr_162  , wr_159  , G207gat );
  not  g202( wr_48   ,           wr_47   );
  nor  g203( wr_174  , wr_173  , wr_170  );
  nor  g204( wr_182  , wr_181  , wr_179  );
  nor  g205( wr_191  , wr_190  , wr_188  );
  nor  g206( wr_201  , wr_200  , wr_199  );
  nor  g207( wr_392  , wr_391  , wr_41   );
  nor  g208( wr_430  , wr_388  , wr_177  );
  nor  g209( wr_403  , wr_388  , wr_275  );
  nor  g210( wr_413  , wr_388  , wr_283  );
  nor  g211( wr_389  , wr_388  , wr_254  );
  nor  g212( wr_237  , wr_236  , wr_71   );
  nor  g213( wr_98   , wr_97   , wr_81   );
  nor  g214( wr_118  , wr_117  , wr_101  );
  nor  g215( wr_141  , wr_140  , wr_81   );
  nor  g216( wr_161  , wr_160  , wr_144  );
  nor  g217( wr_49   , wr_48   , G390gat );
  nor  g218( wr_61   , wr_48   , wr_60   );
  nor  g219( G448gat , wr_74   , wr_71   );
  nor  g220( G449gat , wr_79   , wr_71   );
  not  g221( wr_175  ,           wr_174  );
  nor  g222( wr_183  , wr_182  , wr_39   );
  not  g223( wr_192  ,           wr_191  );
  not  g224( wr_393  ,           wr_392  );
  not  g225( wr_238  ,           wr_237  );
  nor  g226( wr_100  , wr_99   , wr_98   );
  nor  g227( wr_120  , wr_119  , wr_118  );
  nor  g228( wr_143  , wr_142  , wr_141  );
  nor  g229( wr_163  , wr_162  , wr_161  );
  not  g230( G419gat ,           wr_49   );
  not  g231( G446gat ,           wr_61   );
  nor  g232( wr_176  , wr_175  , G268gat );
  nor  g233( wr_184  , wr_183  , wr_177  );
  nor  g234( wr_193  , wr_192  , wr_50   );
  nor  g235( wr_255  , wr_183  , wr_254  );
  nor  g236( wr_276  , wr_183  , wr_275  );
  nor  g237( wr_284  , wr_183  , wr_283  );
  nor  g238( wr_394  , wr_393  , G268gat );
  nor  g239( wr_239  , wr_238  , wr_229  );
  not  g240( wr_122  ,           wr_100  );
  not  g241( wr_123  ,           wr_120  );
  not  g242( wr_165  ,           wr_143  );
  not  g243( wr_166  ,           wr_163  );
  nor  g244( wr_121  , wr_120  , wr_100  );
  nor  g245( wr_164  , wr_163  , wr_143  );
  nor  g246( wr_202  , wr_201  , wr_193  );
  nor  g247( wr_431  , wr_430  , wr_394  );
  nor  g248( wr_404  , wr_403  , wr_394  );
  nor  g249( wr_414  , wr_413  , wr_394  );
  nor  g250( wr_395  , wr_394  , wr_389  );
  not  g251( wr_240  ,           wr_239  );
  nor  g252( wr_124  , wr_123  , wr_122  );
  nor  g253( wr_167  , wr_166  , wr_165  );
  nor  g254( wr_203  , wr_202  , wr_108  );
  nor  g255( wr_256  , wr_202  , wr_102  );
  nor  g256( wr_277  , wr_202  , wr_103  );
  nor  g257( wr_285  , wr_202  , wr_107  );
  nor  g258( wr_427  , wr_202  , wr_88   );
  nor  g259( wr_400  , wr_202  , wr_83   );
  not  g260( wr_432  ,           wr_431  );
  not  g261( wr_405  ,           wr_404  );
  nor  g262( wr_410  , wr_202  , wr_87   );
  not  g263( wr_415  ,           wr_414  );
  nor  g264( wr_382  , wr_202  , wr_82   );
  not  g265( wr_396  ,           wr_395  );
  nor  g266( wr_241  , wr_240  , wr_151  );
  nor  g267( wr_271  , wr_240  , wr_145  );
  nor  g268( wr_342  , wr_240  , wr_146  );
  nor  g269( wr_369  , wr_240  , wr_150  );
  nor  g270( wr_462  , wr_240  , wr_131  );
  nor  g271( wr_485  , wr_240  , wr_125  );
  nor  g272( wr_509  , wr_240  , wr_126  );
  nor  g273( wr_538  , wr_240  , wr_130  );
  nor  g274( G767gat , wr_124  , wr_121  );
  nor  g275( G768gat , wr_167  , wr_164  );
  nor  g276( wr_204  , wr_203  , wr_184  );
  nor  g277( wr_278  , wr_277  , wr_276  );
  nor  g278( wr_286  , wr_285  , wr_284  );
  nor  g279( wr_257  , wr_256  , wr_255  );
  nor  g280( wr_428  , wr_427  , wr_426  );
  nor  g281( wr_401  , wr_400  , wr_399  );
  nor  g282( wr_411  , wr_410  , wr_409  );
  nor  g283( wr_383  , wr_382  , wr_381  );
  not  g284( wr_205  ,           wr_204  );
  not  g285( wr_279  ,           wr_278  );
  not  g286( wr_287  ,           wr_286  );
  not  g287( wr_258  ,           wr_257  );
  not  g288( wr_429  ,           wr_428  );
  not  g289( wr_402  ,           wr_401  );
  not  g290( wr_412  ,           wr_411  );
  not  g291( wr_384  ,           wr_383  );
  nor  g292( wr_206  , wr_205  , wr_176  );
  nor  g293( wr_280  , wr_279  , wr_176  );
  nor  g294( wr_288  , wr_287  , wr_176  );
  nor  g295( wr_259  , wr_258  , wr_176  );
  nor  g296( wr_433  , wr_432  , wr_429  );
  nor  g297( wr_406  , wr_405  , wr_402  );
  nor  g298( wr_416  , wr_415  , wr_412  );
  nor  g299( wr_397  , wr_396  , wr_384  );
  nor  g300( wr_209  , wr_206  , wr_151  );
  not  g301( wr_281  ,           wr_280  );
  not  g302( wr_207  ,           wr_206  );
  nor  g303( wr_289  , wr_288  , wr_150  );
  nor  g304( wr_292  , wr_280  , wr_146  );
  not  g305( wr_293  ,           wr_288  );
  not  g306( wr_260  ,           wr_259  );
  nor  g307( wr_262  , wr_259  , wr_145  );
  not  g308( wr_434  ,           wr_433  );
  not  g309( wr_407  ,           wr_406  );
  nor  g310( wr_441  , wr_433  , wr_131  );
  not  g311( wr_421  ,           wr_416  );
  nor  g312( wr_417  , wr_416  , wr_130  );
  nor  g313( wr_420  , wr_406  , wr_126  );
  not  g314( wr_451  ,           wr_397  );
  nor  g315( wr_398  , wr_397  , wr_125  );
  nor  g316( wr_246  , wr_206  , wr_245  );
  nor  g317( wr_345  , wr_280  , wr_245  );
  nor  g318( wr_372  , wr_288  , wr_245  );
  nor  g319( wr_270  , wr_259  , wr_245  );
  nor  g320( wr_461  , wr_433  , wr_245  );
  nor  g321( wr_484  , wr_397  , wr_245  );
  nor  g322( wr_508  , wr_406  , wr_245  );
  nor  g323( wr_537  , wr_416  , wr_245  );
  nor  g324( wr_208  , wr_207  , G201gat );
  nor  g325( wr_294  , wr_293  , G195gat );
  not  g326( wr_214  ,           wr_209  );
  nor  g327( wr_282  , wr_281  , G189gat );
  not  g328( wr_290  ,           wr_289  );
  nor  g329( wr_261  , wr_260  , G183gat );
  nor  g330( wr_435  , wr_434  , G177gat );
  nor  g331( wr_408  , wr_407  , G165gat );
  not  g332( wr_442  ,           wr_441  );
  nor  g333( wr_422  , wr_421  , G171gat );
  not  g334( wr_418  ,           wr_417  );
  nor  g335( wr_452  , wr_451  , G159gat );
  nor  g336( wr_247  , wr_246  , wr_244  );
  nor  g337( wr_346  , wr_345  , wr_344  );
  nor  g338( wr_373  , wr_372  , wr_371  );
  not  g339( wr_266  ,           wr_262  );
  nor  g340( wr_272  , wr_271  , wr_270  );
  not  g341( wr_322  ,           wr_292  );
  nor  g342( wr_463  , wr_462  , wr_461  );
  not  g343( wr_480  ,           wr_398  );
  nor  g344( wr_486  , wr_485  , wr_484  );
  not  g345( wr_504  ,           wr_420  );
  nor  g346( wr_510  , wr_509  , wr_508  );
  nor  g347( wr_539  , wr_538  , wr_537  );
  nor  g348( wr_295  , wr_208  , wr_222  );
  nor  g349( wr_300  , wr_282  , wr_214  );
  nor  g350( wr_291  , wr_290  , wr_282  );
  nor  g351( wr_443  , wr_442  , wr_408  );
  nor  g352( wr_328  , wr_294  , wr_222  );
  nor  g353( wr_327  , wr_294  , wr_214  );
  nor  g354( wr_419  , wr_418  , wr_408  );
  nor  g355( wr_513  , wr_442  , wr_422  );
  nor  g356( wr_210  , wr_209  , wr_208  );
  nor  g357( wr_263  , wr_262  , wr_261  );
  nor  g358( wr_319  , wr_292  , wr_282  );
  nor  g359( wr_353  , wr_294  , wr_289  );
  nor  g360( wr_455  , wr_441  , wr_435  );
  nor  g361( wr_477  , wr_452  , wr_398  );
  nor  g362( wr_501  , wr_420  , wr_408  );
  nor  g363( wr_531  , wr_422  , wr_417  );
  not  g364( wr_248  ,           wr_247  );
  not  g365( wr_347  ,           wr_346  );
  not  g366( wr_374  ,           wr_373  );
  nor  g367( wr_215  , wr_214  , wr_213  );
  nor  g368( wr_267  , wr_266  , wr_213  );
  not  g369( wr_273  ,           wr_272  );
  nor  g370( wr_323  , wr_322  , wr_213  );
  nor  g371( wr_356  , wr_290  , wr_213  );
  nor  g372( wr_458  , wr_442  , wr_213  );
  not  g373( wr_464  ,           wr_463  );
  nor  g374( wr_481  , wr_480  , wr_213  );
  not  g375( wr_487  ,           wr_486  );
  nor  g376( wr_505  , wr_504  , wr_213  );
  not  g377( wr_511  ,           wr_510  );
  nor  g378( wr_534  , wr_418  , wr_213  );
  not  g379( wr_540  ,           wr_539  );
  not  g380( wr_301  ,           wr_300  );
  not  g381( wr_296  ,           wr_295  );
  not  g382( wr_444  ,           wr_443  );
  not  g383( wr_329  ,           wr_328  );
  nor  g384( wr_360  , wr_295  , wr_209  );
  not  g385( wr_211  ,           wr_210  );
  not  g386( wr_264  ,           wr_263  );
  not  g387( wr_320  ,           wr_319  );
  not  g388( wr_354  ,           wr_353  );
  not  g389( wr_456  ,           wr_455  );
  not  g390( wr_478  ,           wr_477  );
  not  g391( wr_502  ,           wr_501  );
  not  g392( wr_532  ,           wr_531  );
  nor  g393( wr_221  , wr_210  , G261gat );
  nor  g394( wr_249  , wr_248  , wr_241  );
  nor  g395( wr_348  , wr_347  , wr_342  );
  nor  g396( wr_375  , wr_374  , wr_369  );
  nor  g397( wr_302  , wr_301  , wr_294  );
  nor  g398( wr_297  , wr_296  , wr_282  );
  nor  g399( wr_445  , wr_444  , wr_422  );
  nor  g400( wr_330  , wr_329  , wr_208  );
  not  g401( wr_361  ,           wr_360  );
  nor  g402( wr_223  , wr_211  , wr_222  );
  nor  g403( wr_363  , wr_360  , wr_354  );
  nor  g404( wr_212  , wr_211  , wr_168  );
  not  g405( wr_250  ,           wr_249  );
  nor  g406( wr_265  , wr_264  , wr_168  );
  nor  g407( wr_321  , wr_320  , wr_168  );
  not  g408( wr_349  ,           wr_348  );
  nor  g409( wr_355  , wr_354  , wr_168  );
  not  g410( wr_376  ,           wr_375  );
  nor  g411( wr_457  , wr_456  , wr_168  );
  nor  g412( wr_479  , wr_478  , wr_168  );
  nor  g413( wr_503  , wr_502  , wr_168  );
  nor  g414( wr_533  , wr_532  , wr_168  );
  not  g415( wr_298  ,           wr_297  );
  nor  g416( wr_331  , wr_330  , wr_289  );
  nor  g417( wr_362  , wr_361  , wr_353  );
  nor  g418( wr_224  , wr_223  , wr_221  );
  nor  g419( wr_216  , wr_215  , wr_212  );
  nor  g420( wr_268  , wr_267  , wr_265  );
  nor  g421( wr_324  , wr_323  , wr_321  );
  nor  g422( wr_357  , wr_356  , wr_355  );
  nor  g423( wr_459  , wr_458  , wr_457  );
  nor  g424( wr_482  , wr_481  , wr_479  );
  nor  g425( wr_506  , wr_505  , wr_503  );
  nor  g426( wr_535  , wr_534  , wr_533  );
  nor  g427( wr_299  , wr_298  , wr_294  );
  not  g428( wr_332  ,           wr_331  );
  nor  g429( wr_364  , wr_363  , wr_362  );
  not  g430( wr_225  ,           wr_224  );
  not  g431( wr_217  ,           wr_216  );
  not  g432( wr_269  ,           wr_268  );
  not  g433( wr_325  ,           wr_324  );
  not  g434( wr_358  ,           wr_357  );
  not  g435( wr_460  ,           wr_459  );
  not  g436( wr_483  ,           wr_482  );
  not  g437( wr_507  ,           wr_506  );
  not  g438( wr_536  ,           wr_535  );
  nor  g439( wr_303  , wr_302  , wr_299  );
  nor  g440( wr_333  , wr_332  , wr_327  );
  not  g441( wr_365  ,           wr_364  );
  nor  g442( wr_226  , wr_225  , wr_220  );
  not  g443( wr_304  ,           wr_303  );
  not  g444( wr_334  ,           wr_333  );
  nor  g445( wr_336  , wr_333  , wr_320  );
  nor  g446( wr_366  , wr_365  , wr_220  );
  nor  g447( wr_227  , wr_226  , wr_219  );
  nor  g448( wr_305  , wr_304  , wr_292  );
  nor  g449( wr_335  , wr_334  , wr_319  );
  nor  g450( wr_367  , wr_366  , wr_359  );
  not  g451( wr_228  ,           wr_227  );
  not  g452( wr_306  ,           wr_305  );
  nor  g453( wr_337  , wr_336  , wr_335  );
  not  g454( wr_368  ,           wr_367  );
  nor  g455( wr_251  , wr_250  , wr_228  );
  nor  g456( wr_307  , wr_306  , wr_291  );
  not  g457( wr_338  ,           wr_337  );
  nor  g458( wr_377  , wr_376  , wr_368  );
  not  g459( wr_252  ,           wr_251  );
  nor  g460( wr_423  , wr_307  , wr_261  );
  not  g461( wr_308  ,           wr_307  );
  nor  g462( wr_310  , wr_307  , wr_264  );
  nor  g463( wr_339  , wr_338  , wr_220  );
  not  g464( wr_378  ,           wr_377  );
  nor  g465( wr_253  , wr_252  , wr_217  );
  nor  g466( wr_424  , wr_423  , wr_262  );
  nor  g467( wr_309  , wr_308  , wr_263  );
  nor  g468( wr_340  , wr_339  , wr_326  );
  nor  g469( wr_379  , wr_378  , wr_358  );
  not  g470( G850gat ,           wr_253  );
  nor  g471( wr_436  , wr_435  , wr_424  );
  nor  g472( wr_514  , wr_424  , wr_422  );
  not  g473( wr_466  ,           wr_424  );
  nor  g474( wr_468  , wr_456  , wr_424  );
  nor  g475( wr_311  , wr_310  , wr_309  );
  not  g476( wr_341  ,           wr_340  );
  not  g477( G865gat ,           wr_379  );
  not  g478( wr_437  ,           wr_436  );
  not  g479( wr_515  ,           wr_514  );
  nor  g480( wr_542  , wr_441  , wr_436  );
  nor  g481( wr_467  , wr_455  , wr_466  );
  not  g482( wr_312  ,           wr_311  );
  nor  g483( wr_350  , wr_349  , wr_341  );
  nor  g484( wr_438  , wr_437  , wr_408  );
  nor  g485( wr_516  , wr_515  , wr_435  );
  not  g486( wr_543  ,           wr_542  );
  nor  g487( wr_545  , wr_542  , wr_532  );
  nor  g488( wr_469  , wr_468  , wr_467  );
  nor  g489( wr_313  , wr_312  , wr_220  );
  not  g490( wr_351  ,           wr_350  );
  not  g491( wr_439  ,           wr_438  );
  nor  g492( wr_517  , wr_516  , wr_417  );
  nor  g493( wr_544  , wr_543  , wr_531  );
  not  g494( wr_470  ,           wr_469  );
  nor  g495( wr_314  , wr_313  , wr_274  );
  nor  g496( wr_352  , wr_351  , wr_325  );
  nor  g497( wr_440  , wr_439  , wr_422  );
  not  g498( wr_518  ,           wr_517  );
  nor  g499( wr_546  , wr_545  , wr_544  );
  nor  g500( wr_471  , wr_470  , wr_220  );
  not  g501( wr_315  ,           wr_314  );
  not  g502( G864gat ,           wr_352  );
  nor  g503( wr_446  , wr_445  , wr_440  );
  nor  g504( wr_519  , wr_518  , wr_513  );
  not  g505( wr_547  ,           wr_546  );
  nor  g506( wr_472  , wr_471  , wr_465  );
  nor  g507( wr_316  , wr_315  , wr_273  );
  not  g508( wr_447  ,           wr_446  );
  not  g509( wr_520  ,           wr_519  );
  nor  g510( wr_522  , wr_519  , wr_502  );
  nor  g511( wr_548  , wr_547  , wr_220  );
  not  g512( wr_473  ,           wr_472  );
  not  g513( wr_317  ,           wr_316  );
  nor  g514( wr_448  , wr_447  , wr_420  );
  nor  g515( wr_521  , wr_520  , wr_501  );
  nor  g516( wr_549  , wr_548  , wr_541  );
  nor  g517( wr_474  , wr_473  , wr_464  );
  nor  g518( wr_318  , wr_317  , wr_269  );
  not  g519( wr_449  ,           wr_448  );
  nor  g520( wr_523  , wr_522  , wr_521  );
  not  g521( wr_550  ,           wr_549  );
  not  g522( wr_475  ,           wr_474  );
  not  g523( G863gat ,           wr_318  );
  nor  g524( wr_450  , wr_449  , wr_419  );
  not  g525( wr_524  ,           wr_523  );
  nor  g526( wr_551  , wr_550  , wr_540  );
  nor  g527( wr_476  , wr_475  , wr_460  );
  not  g528( wr_490  ,           wr_450  );
  nor  g529( wr_492  , wr_478  , wr_450  );
  nor  g530( wr_525  , wr_524  , wr_220  );
  nor  g531( wr_453  , wr_452  , wr_450  );
  not  g532( wr_552  ,           wr_551  );
  not  g533( G874gat ,           wr_476  );
  nor  g534( wr_491  , wr_477  , wr_490  );
  nor  g535( wr_526  , wr_525  , wr_512  );
  nor  g536( wr_454  , wr_453  , wr_398  );
  nor  g537( wr_553  , wr_552  , wr_536  );
  nor  g538( wr_493  , wr_492  , wr_491  );
  not  g539( wr_527  ,           wr_526  );
  not  g540( G866gat ,           wr_454  );
  not  g541( G880gat ,           wr_553  );
  not  g542( wr_494  ,           wr_493  );
  nor  g543( wr_528  , wr_527  , wr_511  );
  nor  g544( wr_495  , wr_494  , wr_220  );
  not  g545( wr_529  ,           wr_528  );
  nor  g546( wr_496  , wr_495  , wr_489  );
  nor  g547( wr_530  , wr_529  , wr_507  );
  not  g548( wr_497  ,           wr_496  );
  not  g549( G879gat ,           wr_530  );
  nor  g550( wr_498  , wr_497  , wr_487  );
  not  g551( wr_499  ,           wr_498  );
  nor  g552( wr_500  , wr_499  , wr_483  );
  not  g553( G878gat ,           wr_500  );

endmodule
