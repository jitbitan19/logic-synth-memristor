// NOR_NOT mapped module c7552

module c7552 (
  input  G1      ,
  input  G5      ,
  input  G9      ,
  input  G12     ,
  input  G15     ,
  input  G18     ,
  input  G23     ,
  input  G26     ,
  input  G29     ,
  input  G32     ,
  input  G35     ,
  input  G38     ,
  input  G41     ,
  input  G44     ,
  input  G47     ,
  input  G50     ,
  input  G53     ,
  input  G54     ,
  input  G55     ,
  input  G56     ,
  input  G57     ,
  input  G58     ,
  input  G59     ,
  input  G60     ,
  input  G61     ,
  input  G62     ,
  input  G63     ,
  input  G64     ,
  input  G65     ,
  input  G66     ,
  input  G69     ,
  input  G70     ,
  input  G73     ,
  input  G74     ,
  input  G75     ,
  input  G76     ,
  input  G77     ,
  input  G78     ,
  input  G79     ,
  input  G80     ,
  input  G81     ,
  input  G82     ,
  input  G83     ,
  input  G84     ,
  input  G85     ,
  input  G86     ,
  input  G87     ,
  input  G88     ,
  input  G89     ,
  input  G94     ,
  input  G97     ,
  input  G100    ,
  input  G103    ,
  input  G106    ,
  input  G109    ,
  input  G110    ,
  input  G111    ,
  input  G112    ,
  input  G113    ,
  input  G114    ,
  input  G115    ,
  input  G118    ,
  input  G121    ,
  input  G124    ,
  input  G127    ,
  input  G130    ,
  input  G133    ,
  input  G134    ,
  input  G135    ,
  input  G138    ,
  input  G141    ,
  input  G144    ,
  input  G147    ,
  input  G150    ,
  input  G151    ,
  input  G152    ,
  input  G153    ,
  input  G154    ,
  input  G155    ,
  input  G156    ,
  input  G157    ,
  input  G158    ,
  input  G159    ,
  input  G160    ,
  input  G161    ,
  input  G162    ,
  input  G163    ,
  input  G164    ,
  input  G165    ,
  input  G166    ,
  input  G167    ,
  input  G168    ,
  input  G169    ,
  input  G170    ,
  input  G171    ,
  input  G172    ,
  input  G173    ,
  input  G174    ,
  input  G175    ,
  input  G176    ,
  input  G177    ,
  input  G178    ,
  input  G179    ,
  input  G180    ,
  input  G181    ,
  input  G182    ,
  input  G183    ,
  input  G184    ,
  input  G185    ,
  input  G186    ,
  input  G187    ,
  input  G188    ,
  input  G189    ,
  input  G190    ,
  input  G191    ,
  input  G192    ,
  input  G193    ,
  input  G194    ,
  input  G195    ,
  input  G196    ,
  input  G197    ,
  input  G198    ,
  input  G199    ,
  input  G200    ,
  input  G201    ,
  input  G202    ,
  input  G203    ,
  input  G204    ,
  input  G205    ,
  input  G206    ,
  input  G207    ,
  input  G208    ,
  input  G209    ,
  input  G210    ,
  input  G211    ,
  input  G212    ,
  input  G213    ,
  input  G214    ,
  input  G215    ,
  input  G216    ,
  input  G217    ,
  input  G218    ,
  input  G219    ,
  input  G220    ,
  input  G221    ,
  input  G222    ,
  input  G223    ,
  input  G224    ,
  input  G225    ,
  input  G226    ,
  input  G227    ,
  input  G228    ,
  input  G229    ,
  input  G230    ,
  input  G231    ,
  input  G232    ,
  input  G233    ,
  input  G234    ,
  input  G235    ,
  input  G236    ,
  input  G237    ,
  input  G238    ,
  input  G239    ,
  input  G240    ,
  input  G339    ,
  input  G1197   ,
  input  G1455   ,
  input  G1459   ,
  input  G1462   ,
  input  G1469   ,
  input  G1480   ,
  input  G1486   ,
  input  G1492   ,
  input  G1496   ,
  input  G2204   ,
  input  G2208   ,
  input  G2211   ,
  input  G2218   ,
  input  G2224   ,
  input  G2230   ,
  input  G2236   ,
  input  G2239   ,
  input  G2247   ,
  input  G2253   ,
  input  G2256   ,
  input  G3698   ,
  input  G3701   ,
  input  G3705   ,
  input  G3711   ,
  input  G3717   ,
  input  G3723   ,
  input  G3729   ,
  input  G3737   ,
  input  G3743   ,
  input  G3749   ,
  input  G4393   ,
  input  G4394   ,
  input  G4400   ,
  input  G4405   ,
  input  G4410   ,
  input  G4415   ,
  input  G4420   ,
  input  G4427   ,
  input  G4432   ,
  input  G4437   ,
  input  G4526   ,
  input  G4528   ,
  output G2      ,
  output G3      ,
  output G450    ,
  output G448    ,
  output G444    ,
  output G442    ,
  output G440    ,
  output G438    ,
  output G496    ,
  output G494    ,
  output G492    ,
  output G490    ,
  output G488    ,
  output G486    ,
  output G484    ,
  output G482    ,
  output G480    ,
  output G560    ,
  output G542    ,
  output G558    ,
  output G556    ,
  output G554    ,
  output G552    ,
  output G550    ,
  output G548    ,
  output G546    ,
  output G544    ,
  output G540    ,
  output G538    ,
  output G536    ,
  output G534    ,
  output G532    ,
  output G530    ,
  output G528    ,
  output G526    ,
  output G524    ,
  output G279    ,
  output G436    ,
  output G478    ,
  output G522    ,
  output G402    ,
  output G404    ,
  output G406    ,
  output G408    ,
  output G410    ,
  output G432    ,
  output G446    ,
  output G284    ,
  output G286    ,
  output G289    ,
  output G292    ,
  output G341    ,
  output G281    ,
  output G453    ,
  output G278    ,
  output G373    ,
  output G246    ,
  output G258    ,
  output G264    ,
  output G270    ,
  output G388    ,
  output G391    ,
  output G394    ,
  output G397    ,
  output G376    ,
  output G379    ,
  output G382    ,
  output G385    ,
  output G412    ,
  output G414    ,
  output G416    ,
  output G249    ,
  output G295    ,
  output G324    ,
  output G252    ,
  output G276    ,
  output G310    ,
  output G313    ,
  output G316    ,
  output G319    ,
  output G327    ,
  output G330    ,
  output G333    ,
  output G336    ,
  output G418    ,
  output G273    ,
  output G298    ,
  output G301    ,
  output G304    ,
  output G307    ,
  output G344    ,
  output G422    ,
  output G469    ,
  output G419    ,
  output G471    ,
  output G359    ,
  output G362    ,
  output G365    ,
  output G368    ,
  output G347    ,
  output G350    ,
  output G353    ,
  output G356    ,
  output G321    ,
  output G338    ,
  output G370    ,
  output G399    );

  wire wr_108;
  wire wr_109;
  wire wr_110;
  wire wr_111;
  wire wr_112;
  wire wr_113;
  wire wr_114;
  wire wr_115;
  wire wr_116;
  wire wr_117;
  wire wr_118;
  wire wr_119;
  wire wr_120;
  wire wr_121;
  wire wr_122;
  wire wr_123;
  wire wr_124;
  wire wr_125;
  wire wr_126;
  wire wr_127;
  wire wr_128;
  wire wr_129;
  wire wr_130;
  wire wr_131;
  wire wr_132;
  wire wr_133;
  wire wr_134;
  wire wr_135;
  wire wr_136;
  wire wr_137;
  wire wr_138;
  wire wr_139;
  wire wr_140;
  wire wr_141;
  wire wr_142;
  wire wr_143;
  wire wr_144;
  wire wr_145;
  wire wr_146;
  wire wr_147;
  wire wr_148;
  wire wr_149;
  wire wr_150;
  wire wr_151;
  wire wr_152;
  wire wr_153;
  wire wr_154;
  wire wr_155;
  wire wr_156;
  wire wr_157;
  wire wr_158;
  wire wr_159;
  wire wr_160;
  wire wr_161;
  wire wr_162;
  wire wr_163;
  wire wr_164;
  wire wr_165;
  wire wr_166;
  wire wr_167;
  wire wr_168;
  wire wr_169;
  wire wr_170;
  wire wr_171;
  wire wr_172;
  wire wr_173;
  wire wr_174;
  wire wr_175;
  wire wr_176;
  wire wr_177;
  wire wr_178;
  wire wr_179;
  wire wr_180;
  wire wr_181;
  wire wr_182;
  wire wr_183;
  wire wr_184;
  wire wr_185;
  wire wr_186;
  wire wr_187;
  wire wr_188;
  wire wr_189;
  wire wr_190;
  wire wr_191;
  wire wr_192;
  wire wr_193;
  wire wr_194;
  wire wr_195;
  wire wr_196;
  wire wr_197;
  wire wr_198;
  wire wr_199;
  wire wr_200;
  wire wr_201;
  wire wr_202;
  wire wr_203;
  wire wr_204;
  wire wr_205;
  wire wr_206;
  wire wr_207;
  wire wr_208;
  wire wr_209;
  wire wr_210;
  wire wr_211;
  wire wr_212;
  wire wr_213;
  wire wr_214;
  wire wr_215;
  wire wr_216;
  wire wr_217;
  wire wr_218;
  wire wr_219;
  wire wr_220;
  wire wr_221;
  wire wr_222;
  wire wr_223;
  wire wr_224;
  wire wr_225;
  wire wr_226;
  wire wr_227;
  wire wr_228;
  wire wr_229;
  wire wr_230;
  wire wr_231;
  wire wr_232;
  wire wr_233;
  wire wr_234;
  wire wr_235;
  wire wr_236;
  wire wr_237;
  wire wr_238;
  wire wr_239;
  wire wr_240;
  wire wr_241;
  wire wr_242;
  wire wr_243;
  wire wr_244;
  wire wr_245;
  wire wr_246;
  wire wr_247;
  wire wr_248;
  wire wr_249;
  wire wr_250;
  wire wr_251;
  wire wr_252;
  wire wr_253;
  wire wr_254;
  wire wr_255;
  wire wr_256;
  wire wr_257;
  wire wr_258;
  wire wr_259;
  wire wr_260;
  wire wr_261;
  wire wr_262;
  wire wr_263;
  wire wr_264;
  wire wr_265;
  wire wr_266;
  wire wr_267;
  wire wr_268;
  wire wr_269;
  wire wr_270;
  wire wr_271;
  wire wr_272;
  wire wr_273;
  wire wr_274;
  wire wr_275;
  wire wr_276;
  wire wr_277;
  wire wr_278;
  wire wr_279;
  wire wr_280;
  wire wr_281;
  wire wr_282;
  wire wr_283;
  wire wr_284;
  wire wr_285;
  wire wr_286;
  wire wr_287;
  wire wr_288;
  wire wr_289;
  wire wr_290;
  wire wr_291;
  wire wr_292;
  wire wr_293;
  wire wr_294;
  wire wr_295;
  wire wr_296;
  wire wr_297;
  wire wr_298;
  wire wr_299;
  wire wr_300;
  wire wr_301;
  wire wr_302;
  wire wr_303;
  wire wr_304;
  wire wr_305;
  wire wr_306;
  wire wr_307;
  wire wr_308;
  wire wr_309;
  wire wr_310;
  wire wr_311;
  wire wr_312;
  wire wr_313;
  wire wr_314;
  wire wr_315;
  wire wr_316;
  wire wr_317;
  wire wr_318;
  wire wr_319;
  wire wr_320;
  wire wr_321;
  wire wr_322;
  wire wr_323;
  wire wr_324;
  wire wr_325;
  wire wr_326;
  wire wr_327;
  wire wr_328;
  wire wr_329;
  wire wr_330;
  wire wr_331;
  wire wr_332;
  wire wr_333;
  wire wr_334;
  wire wr_335;
  wire wr_336;
  wire wr_337;
  wire wr_338;
  wire wr_339;
  wire wr_340;
  wire wr_341;
  wire wr_342;
  wire wr_343;
  wire wr_344;
  wire wr_345;
  wire wr_346;
  wire wr_347;
  wire wr_348;
  wire wr_349;
  wire wr_350;
  wire wr_351;
  wire wr_352;
  wire wr_353;
  wire wr_354;
  wire wr_355;
  wire wr_356;
  wire wr_357;
  wire wr_358;
  wire wr_359;
  wire wr_360;
  wire wr_361;
  wire wr_362;
  wire wr_363;
  wire wr_364;
  wire wr_365;
  wire wr_366;
  wire wr_367;
  wire wr_368;
  wire wr_369;
  wire wr_370;
  wire wr_371;
  wire wr_372;
  wire wr_373;
  wire wr_374;
  wire wr_375;
  wire wr_376;
  wire wr_377;
  wire wr_378;
  wire wr_379;
  wire wr_380;
  wire wr_381;
  wire wr_382;
  wire wr_383;
  wire wr_384;
  wire wr_385;
  wire wr_386;
  wire wr_387;
  wire wr_388;
  wire wr_389;
  wire wr_390;
  wire wr_391;
  wire wr_392;
  wire wr_393;
  wire wr_394;
  wire wr_395;
  wire wr_396;
  wire wr_397;
  wire wr_398;
  wire wr_399;
  wire wr_400;
  wire wr_401;
  wire wr_402;
  wire wr_403;
  wire wr_404;
  wire wr_405;
  wire wr_406;
  wire wr_407;
  wire wr_408;
  wire wr_409;
  wire wr_410;
  wire wr_411;
  wire wr_412;
  wire wr_413;
  wire wr_414;
  wire wr_415;
  wire wr_416;
  wire wr_417;
  wire wr_418;
  wire wr_419;
  wire wr_420;
  wire wr_421;
  wire wr_422;
  wire wr_423;
  wire wr_424;
  wire wr_425;
  wire wr_426;
  wire wr_427;
  wire wr_428;
  wire wr_429;
  wire wr_430;
  wire wr_431;
  wire wr_432;
  wire wr_433;
  wire wr_434;
  wire wr_435;
  wire wr_436;
  wire wr_437;
  wire wr_438;
  wire wr_439;
  wire wr_440;
  wire wr_441;
  wire wr_442;
  wire wr_443;
  wire wr_444;
  wire wr_445;
  wire wr_446;
  wire wr_447;
  wire wr_448;
  wire wr_449;
  wire wr_450;
  wire wr_451;
  wire wr_452;
  wire wr_453;
  wire wr_454;
  wire wr_455;
  wire wr_456;
  wire wr_457;
  wire wr_458;
  wire wr_459;
  wire wr_460;
  wire wr_461;
  wire wr_462;
  wire wr_463;
  wire wr_464;
  wire wr_465;
  wire wr_466;
  wire wr_467;
  wire wr_468;
  wire wr_469;
  wire wr_470;
  wire wr_471;
  wire wr_472;
  wire wr_473;
  wire wr_474;
  wire wr_475;
  wire wr_476;
  wire wr_477;
  wire wr_478;
  wire wr_479;
  wire wr_480;
  wire wr_481;
  wire wr_482;
  wire wr_483;
  wire wr_484;
  wire wr_485;
  wire wr_486;
  wire wr_487;
  wire wr_488;
  wire wr_489;
  wire wr_490;
  wire wr_491;
  wire wr_492;
  wire wr_493;
  wire wr_494;
  wire wr_495;
  wire wr_496;
  wire wr_497;
  wire wr_498;
  wire wr_499;
  wire wr_500;
  wire wr_501;
  wire wr_502;
  wire wr_503;
  wire wr_504;
  wire wr_505;
  wire wr_506;
  wire wr_507;
  wire wr_508;
  wire wr_509;
  wire wr_510;
  wire wr_511;
  wire wr_512;
  wire wr_513;
  wire wr_514;
  wire wr_515;
  wire wr_516;
  wire wr_517;
  wire wr_518;
  wire wr_519;
  wire wr_520;
  wire wr_521;
  wire wr_522;
  wire wr_523;
  wire wr_524;
  wire wr_525;
  wire wr_526;
  wire wr_527;
  wire wr_528;
  wire wr_529;
  wire wr_530;
  wire wr_531;
  wire wr_532;
  wire wr_533;
  wire wr_534;
  wire wr_535;
  wire wr_536;
  wire wr_537;
  wire wr_538;
  wire wr_539;
  wire wr_540;
  wire wr_541;
  wire wr_542;
  wire wr_543;
  wire wr_544;
  wire wr_545;
  wire wr_546;
  wire wr_547;
  wire wr_548;
  wire wr_549;
  wire wr_550;
  wire wr_551;
  wire wr_552;
  wire wr_553;
  wire wr_554;
  wire wr_555;
  wire wr_556;
  wire wr_557;
  wire wr_558;
  wire wr_559;
  wire wr_560;
  wire wr_561;
  wire wr_562;
  wire wr_563;
  wire wr_564;
  wire wr_565;
  wire wr_566;
  wire wr_567;
  wire wr_568;
  wire wr_569;
  wire wr_570;
  wire wr_571;
  wire wr_572;
  wire wr_573;
  wire wr_574;
  wire wr_575;
  wire wr_576;
  wire wr_577;
  wire wr_578;
  wire wr_579;
  wire wr_580;
  wire wr_581;
  wire wr_582;
  wire wr_583;
  wire wr_584;
  wire wr_585;
  wire wr_586;
  wire wr_587;
  wire wr_588;
  wire wr_589;
  wire wr_590;
  wire wr_591;
  wire wr_592;
  wire wr_593;
  wire wr_594;
  wire wr_595;
  wire wr_596;
  wire wr_597;
  wire wr_598;
  wire wr_599;
  wire wr_600;
  wire wr_601;
  wire wr_602;
  wire wr_603;
  wire wr_604;
  wire wr_605;
  wire wr_606;
  wire wr_607;
  wire wr_608;
  wire wr_609;
  wire wr_610;
  wire wr_611;
  wire wr_612;
  wire wr_613;
  wire wr_614;
  wire wr_615;
  wire wr_616;
  wire wr_617;
  wire wr_618;
  wire wr_619;
  wire wr_620;
  wire wr_621;
  wire wr_622;
  wire wr_623;
  wire wr_624;
  wire wr_625;
  wire wr_626;
  wire wr_627;
  wire wr_628;
  wire wr_629;
  wire wr_630;
  wire wr_631;
  wire wr_632;
  wire wr_633;
  wire wr_634;
  wire wr_635;
  wire wr_636;
  wire wr_637;
  wire wr_638;
  wire wr_639;
  wire wr_640;
  wire wr_641;
  wire wr_642;
  wire wr_643;
  wire wr_644;
  wire wr_645;
  wire wr_646;
  wire wr_647;
  wire wr_648;
  wire wr_649;
  wire wr_650;
  wire wr_651;
  wire wr_652;
  wire wr_653;
  wire wr_654;
  wire wr_655;
  wire wr_656;
  wire wr_657;
  wire wr_658;
  wire wr_659;
  wire wr_660;
  wire wr_661;
  wire wr_662;
  wire wr_663;
  wire wr_664;
  wire wr_665;
  wire wr_666;
  wire wr_667;
  wire wr_668;
  wire wr_669;
  wire wr_670;
  wire wr_671;
  wire wr_672;
  wire wr_673;
  wire wr_674;
  wire wr_675;
  wire wr_676;
  wire wr_677;
  wire wr_678;
  wire wr_679;
  wire wr_680;
  wire wr_681;
  wire wr_682;
  wire wr_683;
  wire wr_684;
  wire wr_685;
  wire wr_686;
  wire wr_687;
  wire wr_688;
  wire wr_689;
  wire wr_690;
  wire wr_691;
  wire wr_692;
  wire wr_693;
  wire wr_694;
  wire wr_695;
  wire wr_696;
  wire wr_697;
  wire wr_698;
  wire wr_699;
  wire wr_700;
  wire wr_701;
  wire wr_702;
  wire wr_703;
  wire wr_704;
  wire wr_705;
  wire wr_706;
  wire wr_707;
  wire wr_708;
  wire wr_709;
  wire wr_710;
  wire wr_711;
  wire wr_712;
  wire wr_713;
  wire wr_714;
  wire wr_715;
  wire wr_716;
  wire wr_717;
  wire wr_718;
  wire wr_719;
  wire wr_720;
  wire wr_721;
  wire wr_722;
  wire wr_723;
  wire wr_724;
  wire wr_725;
  wire wr_726;
  wire wr_727;
  wire wr_728;
  wire wr_729;
  wire wr_730;
  wire wr_731;
  wire wr_732;
  wire wr_733;
  wire wr_734;
  wire wr_735;
  wire wr_736;
  wire wr_737;
  wire wr_738;
  wire wr_739;
  wire wr_740;
  wire wr_741;
  wire wr_742;
  wire wr_743;
  wire wr_744;
  wire wr_745;
  wire wr_746;
  wire wr_747;
  wire wr_748;
  wire wr_749;
  wire wr_750;
  wire wr_751;
  wire wr_752;
  wire wr_753;
  wire wr_754;
  wire wr_755;
  wire wr_756;
  wire wr_757;
  wire wr_758;
  wire wr_759;
  wire wr_760;
  wire wr_761;
  wire wr_762;
  wire wr_763;
  wire wr_764;
  wire wr_765;
  wire wr_766;
  wire wr_767;
  wire wr_768;
  wire wr_769;
  wire wr_770;
  wire wr_771;
  wire wr_772;
  wire wr_773;
  wire wr_774;
  wire wr_775;
  wire wr_776;
  wire wr_777;
  wire wr_778;
  wire wr_779;
  wire wr_780;
  wire wr_781;
  wire wr_782;
  wire wr_783;
  wire wr_784;
  wire wr_785;
  wire wr_786;
  wire wr_787;
  wire wr_788;
  wire wr_789;
  wire wr_790;
  wire wr_791;
  wire wr_792;
  wire wr_793;
  wire wr_794;
  wire wr_795;
  wire wr_796;
  wire wr_797;
  wire wr_798;
  wire wr_799;
  wire wr_800;
  wire wr_801;
  wire wr_802;
  wire wr_803;
  wire wr_804;
  wire wr_805;
  wire wr_806;
  wire wr_807;
  wire wr_808;
  wire wr_809;
  wire wr_810;
  wire wr_811;
  wire wr_812;
  wire wr_813;
  wire wr_814;
  wire wr_815;
  wire wr_816;
  wire wr_817;
  wire wr_818;
  wire wr_819;
  wire wr_820;
  wire wr_821;
  wire wr_822;
  wire wr_823;
  wire wr_824;
  wire wr_825;
  wire wr_826;
  wire wr_827;
  wire wr_828;
  wire wr_829;
  wire wr_830;
  wire wr_831;
  wire wr_832;
  wire wr_833;
  wire wr_834;
  wire wr_835;
  wire wr_836;
  wire wr_837;
  wire wr_838;
  wire wr_839;
  wire wr_840;
  wire wr_841;
  wire wr_842;
  wire wr_843;
  wire wr_844;
  wire wr_845;
  wire wr_846;
  wire wr_847;
  wire wr_848;
  wire wr_849;
  wire wr_850;
  wire wr_851;
  wire wr_852;
  wire wr_853;
  wire wr_854;
  wire wr_855;
  wire wr_856;
  wire wr_857;
  wire wr_858;
  wire wr_859;
  wire wr_860;
  wire wr_861;
  wire wr_862;
  wire wr_863;
  wire wr_864;
  wire wr_865;
  wire wr_866;
  wire wr_867;
  wire wr_868;
  wire wr_869;
  wire wr_870;
  wire wr_871;
  wire wr_872;
  wire wr_873;
  wire wr_874;
  wire wr_875;
  wire wr_876;
  wire wr_877;
  wire wr_878;
  wire wr_879;
  wire wr_880;
  wire wr_881;
  wire wr_882;
  wire wr_883;
  wire wr_884;
  wire wr_885;
  wire wr_886;
  wire wr_887;
  wire wr_888;
  wire wr_889;
  wire wr_890;
  wire wr_891;
  wire wr_892;
  wire wr_893;
  wire wr_894;
  wire wr_895;
  wire wr_896;
  wire wr_897;
  wire wr_898;
  wire wr_899;
  wire wr_900;
  wire wr_901;
  wire wr_902;
  wire wr_903;
  wire wr_904;
  wire wr_905;
  wire wr_906;
  wire wr_907;
  wire wr_908;
  wire wr_909;
  wire wr_910;
  wire wr_911;
  wire wr_912;
  wire wr_913;
  wire wr_914;
  wire wr_915;
  wire wr_916;
  wire wr_917;
  wire wr_918;
  wire wr_919;
  wire wr_920;
  wire wr_921;
  wire wr_922;
  wire wr_923;
  wire wr_924;
  wire wr_925;
  wire wr_926;
  wire wr_927;
  wire wr_928;
  wire wr_929;
  wire wr_930;
  wire wr_931;
  wire wr_932;
  wire wr_933;
  wire wr_934;
  wire wr_935;
  wire wr_936;
  wire wr_937;
  wire wr_938;
  wire wr_939;
  wire wr_940;
  wire wr_941;
  wire wr_942;
  wire wr_943;
  wire wr_944;
  wire wr_945;
  wire wr_946;
  wire wr_947;
  wire wr_948;
  wire wr_949;
  wire wr_950;
  wire wr_951;
  wire wr_952;
  wire wr_953;
  wire wr_954;
  wire wr_955;
  wire wr_956;
  wire wr_957;
  wire wr_958;
  wire wr_959;
  wire wr_960;
  wire wr_961;
  wire wr_962;
  wire wr_963;
  wire wr_964;
  wire wr_965;
  wire wr_966;
  wire wr_967;
  wire wr_968;
  wire wr_969;
  wire wr_970;
  wire wr_971;
  wire wr_972;
  wire wr_973;
  wire wr_974;
  wire wr_975;
  wire wr_976;
  wire wr_977;
  wire wr_978;
  wire wr_979;
  wire wr_980;
  wire wr_981;
  wire wr_982;
  wire wr_983;
  wire wr_984;
  wire wr_985;
  wire wr_986;
  wire wr_987;
  wire wr_988;
  wire wr_989;
  wire wr_990;
  wire wr_991;
  wire wr_992;
  wire wr_993;
  wire wr_994;
  wire wr_995;
  wire wr_996;
  wire wr_997;
  wire wr_998;
  wire wr_999;
  wire wr_1000;
  wire wr_1001;
  wire wr_1002;
  wire wr_1003;
  wire wr_1004;
  wire wr_1005;
  wire wr_1006;
  wire wr_1007;
  wire wr_1008;
  wire wr_1009;
  wire wr_1010;
  wire wr_1011;
  wire wr_1012;
  wire wr_1013;
  wire wr_1014;
  wire wr_1015;
  wire wr_1016;
  wire wr_1017;
  wire wr_1018;
  wire wr_1019;
  wire wr_1020;
  wire wr_1021;
  wire wr_1022;
  wire wr_1023;
  wire wr_1024;
  wire wr_1025;
  wire wr_1026;
  wire wr_1027;
  wire wr_1028;
  wire wr_1029;
  wire wr_1030;
  wire wr_1031;
  wire wr_1032;
  wire wr_1033;
  wire wr_1034;
  wire wr_1035;
  wire wr_1036;
  wire wr_1037;
  wire wr_1038;
  wire wr_1039;
  wire wr_1040;
  wire wr_1041;
  wire wr_1042;
  wire wr_1043;
  wire wr_1044;
  wire wr_1045;
  wire wr_1046;
  wire wr_1047;
  wire wr_1048;
  wire wr_1049;
  wire wr_1050;
  wire wr_1051;
  wire wr_1052;
  wire wr_1053;
  wire wr_1054;
  wire wr_1055;
  wire wr_1056;
  wire wr_1057;
  wire wr_1058;
  wire wr_1059;
  wire wr_1060;
  wire wr_1061;
  wire wr_1062;
  wire wr_1063;
  wire wr_1064;
  wire wr_1065;
  wire wr_1066;
  wire wr_1067;
  wire wr_1068;
  wire wr_1069;
  wire wr_1070;
  wire wr_1071;
  wire wr_1072;
  wire wr_1073;
  wire wr_1074;
  wire wr_1075;
  wire wr_1076;
  wire wr_1077;
  wire wr_1078;
  wire wr_1079;
  wire wr_1080;
  wire wr_1081;
  wire wr_1082;
  wire wr_1083;
  wire wr_1084;
  wire wr_1085;
  wire wr_1086;
  wire wr_1087;
  wire wr_1088;
  wire wr_1089;
  wire wr_1090;
  wire wr_1091;
  wire wr_1092;
  wire wr_1093;
  wire wr_1094;
  wire wr_1095;
  wire wr_1096;
  wire wr_1097;
  wire wr_1098;
  wire wr_1099;
  wire wr_1100;
  wire wr_1101;
  wire wr_1102;
  wire wr_1103;
  wire wr_1104;
  wire wr_1105;
  wire wr_1106;
  wire wr_1107;
  wire wr_1108;
  wire wr_1109;
  wire wr_1110;
  wire wr_1111;
  wire wr_1112;
  wire wr_1113;
  wire wr_1114;
  wire wr_1115;
  wire wr_1116;
  wire wr_1117;
  wire wr_1118;
  wire wr_1119;
  wire wr_1120;
  wire wr_1121;
  wire wr_1122;
  wire wr_1123;
  wire wr_1124;
  wire wr_1125;
  wire wr_1126;
  wire wr_1127;
  wire wr_1128;
  wire wr_1129;
  wire wr_1130;
  wire wr_1131;
  wire wr_1132;
  wire wr_1133;
  wire wr_1134;
  wire wr_1135;
  wire wr_1136;
  wire wr_1137;
  wire wr_1138;
  wire wr_1139;
  wire wr_1140;
  wire wr_1141;
  wire wr_1142;
  wire wr_1143;
  wire wr_1144;
  wire wr_1145;
  wire wr_1146;
  wire wr_1147;
  wire wr_1148;
  wire wr_1149;
  wire wr_1150;
  wire wr_1151;
  wire wr_1152;
  wire wr_1153;
  wire wr_1154;
  wire wr_1155;
  wire wr_1156;
  wire wr_1157;
  wire wr_1158;
  wire wr_1159;
  wire wr_1160;
  wire wr_1161;
  wire wr_1162;
  wire wr_1163;
  wire wr_1164;
  wire wr_1165;
  wire wr_1166;
  wire wr_1167;
  wire wr_1168;
  wire wr_1169;
  wire wr_1170;
  wire wr_1171;
  wire wr_1172;
  wire wr_1173;
  wire wr_1174;
  wire wr_1175;
  wire wr_1176;
  wire wr_1177;
  wire wr_1178;
  wire wr_1179;
  wire wr_1180;
  wire wr_1181;
  wire wr_1182;
  wire wr_1183;
  wire wr_1184;
  wire wr_1185;
  wire wr_1186;
  wire wr_1187;
  wire wr_1188;
  wire wr_1189;
  wire wr_1190;
  wire wr_1191;
  wire wr_1192;
  wire wr_1193;
  wire wr_1194;
  wire wr_1195;
  wire wr_1196;
  wire wr_1197;
  wire wr_1198;
  wire wr_1199;
  wire wr_1200;
  wire wr_1201;
  wire wr_1202;
  wire wr_1203;
  wire wr_1204;
  wire wr_1205;
  wire wr_1206;
  wire wr_1207;
  wire wr_1208;
  wire wr_1209;
  wire wr_1210;
  wire wr_1211;
  wire wr_1212;
  wire wr_1213;
  wire wr_1214;
  wire wr_1215;
  wire wr_1216;
  wire wr_1217;
  wire wr_1218;
  wire wr_1219;
  wire wr_1220;
  wire wr_1221;
  wire wr_1222;
  wire wr_1223;
  wire wr_1224;
  wire wr_1225;
  wire wr_1226;
  wire wr_1227;
  wire wr_1228;
  wire wr_1229;
  wire wr_1230;
  wire wr_1231;
  wire wr_1232;
  wire wr_1233;
  wire wr_1234;
  wire wr_1235;
  wire wr_1236;
  wire wr_1237;
  wire wr_1238;
  wire wr_1239;
  wire wr_1240;
  wire wr_1241;
  wire wr_1242;
  wire wr_1243;
  wire wr_1244;
  wire wr_1245;
  wire wr_1246;
  wire wr_1247;
  wire wr_1248;
  wire wr_1249;
  wire wr_1250;
  wire wr_1251;
  wire wr_1252;
  wire wr_1253;
  wire wr_1254;
  wire wr_1255;
  wire wr_1256;
  wire wr_1257;
  wire wr_1258;
  wire wr_1259;
  wire wr_1260;
  wire wr_1261;
  wire wr_1262;
  wire wr_1263;
  wire wr_1264;
  wire wr_1265;
  wire wr_1266;
  wire wr_1267;
  wire wr_1268;
  wire wr_1269;
  wire wr_1270;
  wire wr_1271;
  wire wr_1272;
  wire wr_1273;
  wire wr_1274;
  wire wr_1275;
  wire wr_1276;
  wire wr_1277;
  wire wr_1278;
  wire wr_1279;
  wire wr_1280;
  wire wr_1281;
  wire wr_1282;
  wire wr_1283;
  wire wr_1284;
  wire wr_1285;
  wire wr_1286;
  wire wr_1287;
  wire wr_1288;
  wire wr_1289;
  wire wr_1290;
  wire wr_1291;
  wire wr_1292;
  wire wr_1293;
  wire wr_1294;
  wire wr_1295;
  wire wr_1296;
  wire wr_1297;
  wire wr_1298;
  wire wr_1299;
  wire wr_1300;
  wire wr_1301;
  wire wr_1302;
  wire wr_1303;
  wire wr_1304;
  wire wr_1305;
  wire wr_1306;
  wire wr_1307;
  wire wr_1308;
  wire wr_1309;
  wire wr_1310;
  wire wr_1311;
  wire wr_1312;
  wire wr_1313;
  wire wr_1314;
  wire wr_1315;
  wire wr_1316;
  wire wr_1317;
  wire wr_1318;
  wire wr_1319;
  wire wr_1320;
  wire wr_1321;
  wire wr_1322;
  wire wr_1323;
  wire wr_1324;
  wire wr_1325;
  wire wr_1326;
  wire wr_1327;
  wire wr_1328;
  wire wr_1329;
  wire wr_1330;
  wire wr_1331;
  wire wr_1332;
  wire wr_1333;
  wire wr_1334;
  wire wr_1335;
  wire wr_1336;
  wire wr_1337;
  wire wr_1338;
  wire wr_1339;
  wire wr_1340;
  wire wr_1341;
  wire wr_1342;
  wire wr_1343;
  wire wr_1344;
  wire wr_1345;
  wire wr_1346;
  wire wr_1347;
  wire wr_1348;
  wire wr_1349;
  wire wr_1350;
  wire wr_1351;
  wire wr_1352;
  wire wr_1353;
  wire wr_1354;
  wire wr_1355;
  wire wr_1356;
  wire wr_1357;
  wire wr_1358;
  wire wr_1359;
  wire wr_1360;
  wire wr_1361;
  wire wr_1362;
  wire wr_1363;
  wire wr_1364;
  wire wr_1365;
  wire wr_1366;
  wire wr_1367;
  wire wr_1368;
  wire wr_1369;
  wire wr_1370;
  wire wr_1371;
  wire wr_1372;
  wire wr_1373;
  wire wr_1374;
  wire wr_1375;
  wire wr_1376;
  wire wr_1377;
  wire wr_1378;
  wire wr_1379;
  wire wr_1380;
  wire wr_1381;
  wire wr_1382;
  wire wr_1383;
  wire wr_1384;
  wire wr_1385;
  wire wr_1386;
  wire wr_1387;
  wire wr_1388;
  wire wr_1389;
  wire wr_1390;
  wire wr_1391;
  wire wr_1392;
  wire wr_1393;
  wire wr_1394;
  wire wr_1395;
  wire wr_1396;
  wire wr_1397;
  wire wr_1398;
  wire wr_1399;
  wire wr_1400;
  wire wr_1401;
  wire wr_1402;
  wire wr_1403;
  wire wr_1404;
  wire wr_1405;
  wire wr_1406;
  wire wr_1407;
  wire wr_1408;
  wire wr_1409;
  wire wr_1410;
  wire wr_1411;
  wire wr_1412;
  wire wr_1413;
  wire wr_1414;
  wire wr_1415;
  wire wr_1416;
  wire wr_1417;
  wire wr_1418;
  wire wr_1419;
  wire wr_1420;
  wire wr_1421;
  wire wr_1422;
  wire wr_1423;
  wire wr_1424;
  wire wr_1425;
  wire wr_1426;
  wire wr_1427;
  wire wr_1428;
  wire wr_1429;
  wire wr_1430;
  wire wr_1431;
  wire wr_1432;
  wire wr_1433;
  wire wr_1434;
  wire wr_1435;
  wire wr_1436;
  wire wr_1437;
  wire wr_1438;
  wire wr_1439;
  wire wr_1440;
  wire wr_1441;
  wire wr_1442;
  wire wr_1443;
  wire wr_1444;
  wire wr_1445;
  wire wr_1446;
  wire wr_1447;
  wire wr_1448;
  wire wr_1449;
  wire wr_1450;
  wire wr_1451;
  wire wr_1452;
  wire wr_1453;
  wire wr_1454;
  wire wr_1455;
  wire wr_1456;
  wire wr_1457;
  wire wr_1458;
  wire wr_1459;
  wire wr_1460;
  wire wr_1461;
  wire wr_1462;
  wire wr_1463;
  wire wr_1464;
  wire wr_1465;
  wire wr_1466;
  wire wr_1467;
  wire wr_1468;
  wire wr_1469;
  wire wr_1470;
  wire wr_1471;
  wire wr_1472;
  wire wr_1473;
  wire wr_1474;
  wire wr_1475;
  wire wr_1476;
  wire wr_1477;
  wire wr_1478;
  wire wr_1479;
  wire wr_1480;
  wire wr_1481;
  wire wr_1482;
  wire wr_1483;
  wire wr_1484;
  wire wr_1485;
  wire wr_1486;
  wire wr_1487;
  wire wr_1488;
  wire wr_1489;
  wire wr_1490;
  wire wr_1491;
  wire wr_1492;
  wire wr_1493;
  wire wr_1494;
  wire wr_1495;
  wire wr_1496;
  wire wr_1497;
  wire wr_1498;
  wire wr_1499;
  wire wr_1500;
  wire wr_1501;
  wire wr_1502;
  wire wr_1503;
  wire wr_1504;
  wire wr_1505;
  wire wr_1506;
  wire wr_1507;
  wire wr_1508;
  wire wr_1509;
  wire wr_1510;
  wire wr_1511;
  wire wr_1512;
  wire wr_1513;
  wire wr_1514;
  wire wr_1515;
  wire wr_1516;
  wire wr_1517;
  wire wr_1518;
  wire wr_1519;
  wire wr_1520;
  wire wr_1521;
  wire wr_1522;
  wire wr_1523;
  wire wr_1524;
  wire wr_1525;
  wire wr_1526;
  wire wr_1527;
  wire wr_1528;
  wire wr_1529;
  wire wr_1530;
  wire wr_1531;
  wire wr_1532;
  wire wr_1533;
  wire wr_1534;
  wire wr_1535;
  wire wr_1536;
  wire wr_1537;
  wire wr_1538;
  wire wr_1539;
  wire wr_1540;
  wire wr_1541;
  wire wr_1542;
  wire wr_1543;
  wire wr_1544;
  wire wr_1545;
  wire wr_1546;
  wire wr_1547;
  wire wr_1548;
  wire wr_1549;
  wire wr_1550;
  wire wr_1551;
  wire wr_1552;
  wire wr_1553;
  wire wr_1554;
  wire wr_1555;
  wire wr_1556;
  wire wr_1557;
  wire wr_1558;
  wire wr_1559;
  wire wr_1560;
  wire wr_1561;
  wire wr_1562;
  wire wr_1563;
  wire wr_1564;
  wire wr_1565;
  wire wr_1566;
  wire wr_1567;
  wire wr_1568;
  wire wr_1569;
  wire wr_1570;
  wire wr_1571;
  wire wr_1572;
  wire wr_1573;
  wire wr_1574;
  wire wr_1575;
  wire wr_1576;
  wire wr_1577;
  wire wr_1578;
  wire wr_1579;
  wire wr_1580;
  wire wr_1581;
  wire wr_1582;
  wire wr_1583;
  wire wr_1584;
  wire wr_1585;
  wire wr_1586;
  wire wr_1587;
  wire wr_1588;
  wire wr_1589;
  wire wr_1590;
  wire wr_1591;
  wire wr_1592;
  wire wr_1593;
  wire wr_1594;
  wire wr_1595;
  wire wr_1596;
  wire wr_1597;
  wire wr_1598;
  wire wr_1599;
  wire wr_1600;
  wire wr_1601;
  wire wr_1602;
  wire wr_1603;
  wire wr_1604;
  wire wr_1605;
  wire wr_1606;
  wire wr_1607;
  wire wr_1608;
  wire wr_1609;
  wire wr_1610;
  wire wr_1611;
  wire wr_1612;
  wire wr_1613;
  wire wr_1614;
  wire wr_1615;
  wire wr_1616;
  wire wr_1617;
  wire wr_1618;
  wire wr_1619;
  wire wr_1620;
  wire wr_1621;
  wire wr_1622;
  wire wr_1623;
  wire wr_1624;
  wire wr_1625;
  wire wr_1626;
  wire wr_1627;
  wire wr_1628;
  wire wr_1629;
  wire wr_1630;
  wire wr_1631;
  wire wr_1632;
  wire wr_1633;
  wire wr_1634;
  wire wr_1635;
  wire wr_1636;
  wire wr_1637;
  wire wr_1638;
  wire wr_1639;
  wire wr_1640;
  wire wr_1641;
  wire wr_1642;
  wire wr_1643;
  wire wr_1644;
  wire wr_1645;
  wire wr_1646;
  wire wr_1647;
  wire wr_1648;
  wire wr_1649;
  wire wr_1650;
  wire wr_1651;
  wire wr_1652;
  wire wr_1653;
  wire wr_1654;
  wire wr_1655;
  wire wr_1656;
  wire wr_1657;
  wire wr_1658;
  wire wr_1659;
  wire wr_1660;
  wire wr_1661;
  wire wr_1662;
  wire wr_1663;
  wire wr_1664;
  wire wr_1665;
  wire wr_1666;
  wire wr_1667;
  wire wr_1668;
  wire wr_1669;
  wire wr_1670;
  wire wr_1671;
  wire wr_1672;
  wire wr_1673;
  wire wr_1674;
  wire wr_1675;
  wire wr_1676;
  wire wr_1677;
  wire wr_1678;
  wire wr_1679;
  wire wr_1680;
  wire wr_1681;
  wire wr_1682;
  wire wr_1683;
  wire wr_1684;
  wire wr_1685;
  wire wr_1686;
  wire wr_1687;
  wire wr_1688;
  wire wr_1689;
  wire wr_1690;
  wire wr_1691;
  wire wr_1692;
  wire wr_1693;
  wire wr_1694;
  wire wr_1695;
  wire wr_1696;
  wire wr_1697;
  wire wr_1698;
  wire wr_1699;
  wire wr_1700;
  wire wr_1701;
  wire wr_1702;
  wire wr_1703;
  wire wr_1704;
  wire wr_1705;
  wire wr_1706;
  wire wr_1707;
  wire wr_1708;
  wire wr_1709;
  wire wr_1710;
  wire wr_1711;
  wire wr_1712;
  wire wr_1713;
  wire wr_1714;
  wire wr_1715;
  wire wr_1716;
  wire wr_1717;
  wire wr_1718;
  wire wr_1719;
  wire wr_1720;
  wire wr_1721;
  wire wr_1722;
  wire wr_1723;
  wire wr_1724;
  wire wr_1725;
  wire wr_1726;
  wire wr_1727;
  wire wr_1728;
  wire wr_1729;
  wire wr_1730;
  wire wr_1731;
  wire wr_1732;
  wire wr_1733;
  wire wr_1734;
  wire wr_1735;
  wire wr_1736;
  wire wr_1737;
  wire wr_1738;
  wire wr_1739;
  wire wr_1740;
  wire wr_1741;
  wire wr_1742;
  wire wr_1743;
  wire wr_1744;
  wire wr_1745;
  wire wr_1746;
  wire wr_1747;
  wire wr_1748;
  wire wr_1749;
  wire wr_1750;
  wire wr_1751;
  wire wr_1752;
  wire wr_1753;
  wire wr_1754;
  wire wr_1755;
  wire wr_1756;
  wire wr_1757;
  wire wr_1758;
  wire wr_1759;
  wire wr_1760;
  wire wr_1761;
  wire wr_1762;
  wire wr_1763;
  wire wr_1764;
  wire wr_1765;
  wire wr_1766;
  wire wr_1767;
  wire wr_1768;
  wire wr_1769;
  wire wr_1770;
  wire wr_1771;
  wire wr_1772;
  wire wr_1773;
  wire wr_1774;
  wire wr_1775;
  wire wr_1776;
  wire wr_1777;
  wire wr_1778;
  wire wr_1779;
  wire wr_1780;
  wire wr_1781;
  wire wr_1782;
  wire wr_1783;
  wire wr_1784;
  wire wr_1785;
  wire wr_1786;
  wire wr_1787;
  wire wr_1788;
  wire wr_1789;
  wire wr_1790;
  wire wr_1791;
  wire wr_1792;
  wire wr_1793;
  wire wr_1794;
  wire wr_1795;
  wire wr_1796;
  wire wr_1797;
  wire wr_1798;
  wire wr_1799;
  wire wr_1800;
  wire wr_1801;
  wire wr_1802;
  wire wr_1803;
  wire wr_1804;
  wire wr_1805;
  wire wr_1806;
  wire wr_1807;
  wire wr_1808;
  wire wr_1809;
  wire wr_1810;
  wire wr_1811;
  wire wr_1812;
  wire wr_1813;
  wire wr_1814;
  wire wr_1815;
  wire wr_1816;
  wire wr_1817;
  wire wr_1818;
  wire wr_1819;
  wire wr_1820;
  wire wr_1821;
  wire wr_1822;
  wire wr_1823;
  wire wr_1824;
  wire wr_1825;
  wire wr_1826;
  wire wr_1827;
  wire wr_1828;
  wire wr_1829;
  wire wr_1830;
  wire wr_1831;
  wire wr_1832;
  wire wr_1833;
  wire wr_1834;
  wire wr_1835;
  wire wr_1836;
  wire wr_1837;
  wire wr_1838;
  wire wr_1839;
  wire wr_1840;
  wire wr_1841;
  wire wr_1842;
  wire wr_1843;
  wire wr_1844;
  wire wr_1845;
  wire wr_1846;
  wire wr_1847;
  wire wr_1848;
  wire wr_1849;
  wire wr_1850;
  wire wr_1851;
  wire wr_1852;
  wire wr_1853;
  wire wr_1854;
  wire wr_1855;
  wire wr_1856;
  wire wr_1857;
  wire wr_1858;
  wire wr_1859;
  wire wr_1860;
  wire wr_1861;
  wire wr_1862;
  wire wr_1863;
  wire wr_1864;
  wire wr_1865;
  wire wr_1866;
  wire wr_1867;
  wire wr_1868;
  wire wr_1869;
  wire wr_1870;
  wire wr_1871;
  wire wr_1872;
  wire wr_1873;
  wire wr_1874;
  wire wr_1875;
  wire wr_1876;
  wire wr_1877;
  wire wr_1878;
  wire wr_1879;
  wire wr_1880;
  wire wr_1881;
  wire wr_1882;
  wire wr_1883;
  wire wr_1884;
  wire wr_1885;
  wire wr_1886;
  wire wr_1887;
  wire wr_1888;
  wire wr_1889;
  wire wr_1890;
  wire wr_1891;
  wire wr_1892;
  wire wr_1893;
  wire wr_1894;
  wire wr_1895;
  wire wr_1896;
  wire wr_1897;
  wire wr_1898;
  wire wr_1899;
  wire wr_1900;
  wire wr_1901;
  wire wr_1902;
  wire wr_1903;
  wire wr_1904;
  wire wr_1905;
  wire wr_1906;
  wire wr_1907;
  wire wr_1908;
  wire wr_1909;
  wire wr_1910;
  wire wr_1911;
  wire wr_1912;
  wire wr_1913;
  wire wr_1914;
  wire wr_1915;
  wire wr_1916;
  wire wr_1917;
  wire wr_1918;
  wire wr_1919;
  wire wr_1920;
  wire wr_1921;
  wire wr_1922;
  wire wr_1923;
  wire wr_1924;
  wire wr_1925;
  wire wr_1926;
  wire wr_1927;
  wire wr_1928;
  wire wr_1929;
  wire wr_1930;
  wire wr_1931;
  wire wr_1932;
  wire wr_1933;
  wire wr_1934;
  wire wr_1935;
  wire wr_1936;
  wire wr_1937;
  wire wr_1938;
  wire wr_1939;
  wire wr_1940;
  wire wr_1941;
  wire wr_1942;
  wire wr_1943;
  wire wr_1944;
  wire wr_1945;
  wire wr_1946;
  wire wr_1947;
  wire wr_1948;
  wire wr_1949;
  wire wr_1950;
  wire wr_1951;
  wire wr_1952;
  wire wr_1953;
  wire wr_1954;
  wire wr_1955;
  wire wr_1956;
  wire wr_1957;
  wire wr_1958;
  wire wr_1959;
  wire wr_1960;
  wire wr_1961;
  wire wr_1962;
  wire wr_1963;
  wire wr_1964;
  wire wr_1965;
  wire wr_1966;
  wire wr_1967;
  wire wr_1968;
  wire wr_1969;
  wire wr_1970;
  wire wr_1971;
  wire wr_1972;
  wire wr_1973;
  wire wr_1974;
  wire wr_1975;
  wire wr_1976;
  wire wr_1977;
  wire wr_1978;
  wire wr_1979;
  wire wr_1980;
  wire wr_1981;
  wire wr_1982;
  wire wr_1983;
  wire wr_1984;
  wire wr_1985;
  wire wr_1986;
  wire wr_1987;
  wire wr_1988;
  wire wr_1989;
  wire wr_1990;
  wire wr_1991;
  wire wr_1992;
  wire wr_1993;
  wire wr_1994;
  wire wr_1995;
  wire wr_1996;
  wire wr_1997;
  wire wr_1998;
  wire wr_1999;
  wire wr_2000;
  wire wr_2001;
  wire wr_2002;
  wire wr_2003;
  wire wr_2004;
  wire wr_2005;
  wire wr_2006;
  wire wr_2007;
  wire wr_2008;
  wire wr_2009;
  wire wr_2010;
  wire wr_2011;
  wire wr_2012;
  wire wr_2013;
  wire wr_2014;
  wire wr_2015;
  wire wr_2016;
  wire wr_2017;
  wire wr_2018;
  wire wr_2019;
  wire wr_2020;
  wire wr_2021;
  wire wr_2022;
  wire wr_2023;
  wire wr_2024;
  wire wr_2025;
  wire wr_2026;
  wire wr_2027;
  wire wr_2028;
  wire wr_2029;
  wire wr_2030;
  wire wr_2031;
  wire wr_2032;
  wire wr_2033;
  wire wr_2034;
  wire wr_2035;
  wire wr_2036;
  wire wr_2037;
  wire wr_2038;
  wire wr_2039;
  wire wr_2040;
  wire wr_2041;
  wire wr_2042;
  wire wr_2043;
  wire wr_2044;
  wire wr_2045;
  wire wr_2046;
  wire wr_2047;
  wire wr_2048;
  wire wr_2049;
  wire wr_2050;
  wire wr_2051;
  wire wr_2052;
  wire wr_2053;
  wire wr_2054;
  wire wr_2055;
  wire wr_2056;
  wire wr_2057;
  wire wr_2058;
  wire wr_2059;
  wire wr_2060;
  wire wr_2061;
  wire wr_2062;
  wire wr_2063;
  wire wr_2064;
  wire wr_2065;
  wire wr_2066;
  wire wr_2067;
  wire wr_2068;
  wire wr_2069;
  wire wr_2070;
  wire wr_2071;
  wire wr_2072;
  wire wr_2073;
  wire wr_2074;
  wire wr_2075;
  wire wr_2076;
  wire wr_2077;
  wire wr_2078;
  wire wr_2079;
  wire wr_2080;
  wire wr_2081;
  wire wr_2082;
  wire wr_2083;
  wire wr_2084;
  wire wr_2085;
  wire wr_2086;
  wire wr_2087;
  wire wr_2088;
  wire wr_2089;
  wire wr_2090;
  wire wr_2091;
  wire wr_2092;
  wire wr_2093;
  wire wr_2094;
  wire wr_2095;
  wire wr_2096;
  wire wr_2097;
  wire wr_2098;
  wire wr_2099;
  wire wr_2100;
  wire wr_2101;
  wire wr_2102;
  wire wr_2103;
  wire wr_2104;
  wire wr_2105;
  wire wr_2106;
  wire wr_2107;
  wire wr_2108;
  wire wr_2109;
  wire wr_2110;
  wire wr_2111;
  wire wr_2112;
  wire wr_2113;
  wire wr_2114;
  wire wr_2115;
  wire wr_2116;
  wire wr_2117;
  wire wr_2118;
  wire wr_2119;
  wire wr_2120;
  wire wr_2121;
  wire wr_2122;
  wire wr_2123;
  wire wr_2124;
  wire wr_2125;
  wire wr_2126;
  wire wr_2127;
  wire wr_2128;
  wire wr_2129;
  wire wr_2130;
  wire wr_2131;
  wire wr_2132;
  wire wr_2133;
  wire wr_2134;
  wire wr_2135;
  wire wr_2136;
  wire wr_2137;
  wire wr_2138;
  wire wr_2139;
  wire wr_2140;
  wire wr_2141;
  wire wr_2142;
  wire wr_2143;
  wire wr_2144;
  wire wr_2145;
  wire wr_2146;
  wire wr_2147;
  wire wr_2148;
  wire wr_2149;
  wire wr_2150;
  wire wr_2151;
  wire wr_2152;
  wire wr_2153;
  wire wr_2154;
  wire wr_2155;
  wire wr_2156;
  wire wr_2157;
  wire wr_2158;
  wire wr_2159;
  wire wr_2160;
  wire wr_2161;
  wire wr_2162;
  wire wr_2163;
  wire wr_2164;
  wire wr_2165;
  wire wr_2166;
  wire wr_2167;
  wire wr_2168;
  wire wr_2169;
  wire wr_2170;
  wire wr_2171;
  wire wr_2172;
  wire wr_2173;
  wire wr_2174;
  wire wr_2175;
  wire wr_2176;
  wire wr_2177;
  wire wr_2178;
  wire wr_2179;
  wire wr_2180;
  wire wr_2181;
  wire wr_2182;
  wire wr_2183;
  wire wr_2184;
  wire wr_2185;
  wire wr_2186;
  wire wr_2187;
  wire wr_2188;
  wire wr_2189;
  wire wr_2190;
  wire wr_2191;
  wire wr_2192;
  wire wr_2193;
  wire wr_2194;
  wire wr_2195;
  wire wr_2196;
  wire wr_2197;
  wire wr_2198;
  wire wr_2199;
  wire wr_2200;
  wire wr_2201;
  wire wr_2202;
  wire wr_2203;
  wire wr_2204;
  wire wr_2205;
  wire wr_2206;
  wire wr_2207;
  wire wr_2208;
  wire wr_2209;
  wire wr_2210;
  wire wr_2211;
  wire wr_2212;
  wire wr_2213;
  wire wr_2214;
  wire wr_2215;
  wire wr_2216;
  wire wr_2217;
  wire wr_2218;
  wire wr_2219;
  wire wr_2220;
  wire wr_2221;
  wire wr_2222;
  wire wr_2223;
  wire wr_2224;
  wire wr_2225;
  wire wr_2226;
  wire wr_2227;
  wire wr_2228;
  wire wr_2229;
  wire wr_2230;
  wire wr_2231;
  wire wr_2232;
  wire wr_2233;
  wire wr_2234;
  wire wr_2235;
  wire wr_2236;
  wire wr_2237;
  wire wr_2238;
  wire wr_2239;
  wire wr_2240;
  wire wr_2241;
  wire wr_2242;
  wire wr_2243;
  wire wr_2244;
  wire wr_2245;
  wire wr_2246;
  wire wr_2247;
  wire wr_2248;
  wire wr_2249;
  wire wr_2250;
  wire wr_2251;
  wire wr_2252;
  wire wr_2253;
  wire wr_2254;
  wire wr_2255;
  wire wr_2256;
  wire wr_2257;
  wire wr_2258;
  wire wr_2259;
  wire wr_2260;
  wire wr_2261;
  wire wr_2262;
  wire wr_2263;
  wire wr_2264;
  wire wr_2265;
  wire wr_2266;
  wire wr_2267;
  wire wr_2268;
  wire wr_2269;
  wire wr_2270;
  wire wr_2271;
  wire wr_2272;
  wire wr_2273;
  wire wr_2274;
  wire wr_2275;
  wire wr_2276;
  wire wr_2277;
  wire wr_2278;
  wire wr_2279;
  wire wr_2280;
  wire wr_2281;
  wire wr_2282;
  wire wr_2283;
  wire wr_2284;
  wire wr_2285;
  wire wr_2286;
  wire wr_2287;
  wire wr_2288;
  wire wr_2289;
  wire wr_2290;
  wire wr_2291;
  wire wr_2292;
  wire wr_2293;
  wire wr_2294;
  wire wr_2295;
  wire wr_2296;
  wire wr_2297;
  wire wr_2298;
  wire wr_2299;
  wire wr_2300;
  wire wr_2301;
  wire wr_2302;
  wire wr_2303;
  wire wr_2304;
  wire wr_2305;
  wire wr_2306;
  wire wr_2307;
  wire wr_2308;
  wire wr_2309;
  wire wr_2310;
  wire wr_2311;
  wire wr_2312;
  wire wr_2313;
  wire wr_2314;
  wire wr_2315;
  wire wr_2316;
  wire wr_2317;
  wire wr_2318;
  wire wr_2319;
  wire wr_2320;
  wire wr_2321;
  wire wr_2322;
  wire wr_2323;
  wire wr_2324;
  wire wr_2325;
  wire wr_2326;
  wire wr_2327;
  wire wr_2328;
  wire wr_2329;
  wire wr_2330;
  wire wr_2331;
  wire wr_2332;
  wire wr_2333;
  wire wr_2334;
  wire wr_2335;
  wire wr_2336;
  wire wr_2337;
  wire wr_2338;
  wire wr_2339;
  wire wr_2340;
  wire wr_2341;
  wire wr_2342;
  wire wr_2343;
  wire wr_2344;
  wire wr_2345;
  wire wr_2346;
  wire wr_2347;
  wire wr_2348;
  wire wr_2349;
  wire wr_2350;
  wire wr_2351;
  wire wr_2352;
  wire wr_2353;
  wire wr_2354;
  wire wr_2355;
  wire wr_2356;
  wire wr_2357;
  wire wr_2358;
  wire wr_2359;
  wire wr_2360;
  wire wr_2361;
  wire wr_2362;
  wire wr_2363;
  wire wr_2364;
  wire wr_2365;
  wire wr_2366;
  wire wr_2367;
  wire wr_2368;
  wire wr_2369;
  wire wr_2370;
  wire wr_2371;
  wire wr_2372;
  wire wr_2373;
  wire wr_2374;
  wire wr_2375;
  wire wr_2376;
  wire wr_2377;
  wire wr_2378;
  wire wr_2379;
  wire wr_2380;
  wire wr_2381;
  wire wr_2382;
  wire wr_2383;
  wire wr_2384;
  wire wr_2385;
  wire wr_2386;
  wire wr_2387;
  wire wr_2388;
  wire wr_2389;
  wire wr_2390;
  wire wr_2391;
  wire wr_2392;
  wire wr_2393;
  wire wr_2394;
  wire wr_2395;
  wire wr_2396;
  wire wr_2397;
  wire wr_2398;
  wire wr_2399;
  wire wr_2400;
  wire wr_2401;
  wire wr_2402;
  wire wr_2403;
  wire wr_2404;
  wire wr_2405;
  wire wr_2406;
  wire wr_2407;
  wire wr_2408;
  wire wr_2409;
  wire wr_2410;
  wire wr_2411;
  wire wr_2412;
  wire wr_2413;
  wire wr_2414;
  wire wr_2415;
  wire wr_2416;
  wire wr_2417;
  wire wr_2418;
  wire wr_2419;
  wire wr_2420;
  wire wr_2421;
  wire wr_2422;
  wire wr_2423;
  wire wr_2424;
  wire wr_2425;
  wire wr_2426;
  wire wr_2427;
  wire wr_2428;
  wire wr_2429;
  wire wr_2430;
  wire wr_2431;
  wire wr_2432;
  wire wr_2433;
  wire wr_2434;
  wire wr_2435;
  wire wr_2436;
  wire wr_2437;
  wire wr_2438;
  wire wr_2439;
  wire wr_2440;
  wire wr_2441;
  wire wr_2442;
  wire wr_2443;
  wire wr_2444;
  wire wr_2445;
  wire wr_2446;
  wire wr_2447;
  wire wr_2448;
  wire wr_2449;
  wire wr_2450;
  wire wr_2451;
  wire wr_2452;
  wire wr_2453;
  wire wr_2454;
  wire wr_2455;
  wire wr_2456;
  wire wr_2457;
  wire wr_2458;
  wire wr_2459;
  wire wr_2460;
  wire wr_2461;
  wire wr_2462;
  wire wr_2463;
  wire wr_2464;
  wire wr_2465;
  wire wr_2466;
  wire wr_2467;
  wire wr_2468;
  wire wr_2469;
  wire wr_2470;
  wire wr_2471;
  wire wr_2472;
  wire wr_2473;
  wire wr_2474;
  wire wr_2475;
  wire wr_2476;
  wire wr_2477;
  wire wr_2478;
  wire wr_2479;
  wire wr_2480;
  wire wr_2481;
  wire wr_2482;
  wire wr_2483;
  wire wr_2484;
  wire wr_2485;
  wire wr_2486;
  wire wr_2487;
  wire wr_2488;
  wire wr_2489;
  wire wr_2490;
  wire wr_2491;
  wire wr_2492;
  wire wr_2493;
  wire wr_2494;
  wire wr_2495;
  wire wr_2496;
  wire wr_2497;
  wire wr_2498;
  wire wr_2499;
  wire wr_2500;
  wire wr_2501;
  wire wr_2502;
  wire wr_2503;
  wire wr_2504;
  wire wr_2505;
  wire wr_2506;
  wire wr_2507;
  wire wr_2508;
  wire wr_2509;
  wire wr_2510;
  wire wr_2511;
  wire wr_2512;
  wire wr_2513;
  wire wr_2514;
  wire wr_2515;
  wire wr_2516;
  wire wr_2517;
  wire wr_2518;
  wire wr_2519;
  wire wr_2520;
  wire wr_2521;
  wire wr_2522;
  wire wr_2523;
  wire wr_2524;
  wire wr_2525;
  wire wr_2526;
  wire wr_2527;
  wire wr_2528;
  wire wr_2529;
  wire wr_2530;
  wire wr_2531;
  wire wr_2532;
  wire wr_2533;
  wire wr_2534;
  wire wr_2535;
  wire wr_2536;
  wire wr_2537;
  wire wr_2538;
  wire wr_2539;
  wire wr_2540;
  wire wr_2541;
  wire wr_2542;
  wire wr_2543;
  wire wr_2544;
  wire wr_2545;
  wire wr_2546;
  wire wr_2547;
  wire wr_2548;
  wire wr_2549;
  wire wr_2550;
  wire wr_2551;
  wire wr_2552;
  wire wr_2553;
  wire wr_2554;
  wire wr_2555;
  wire wr_2556;
  wire wr_2557;
  wire wr_2558;
  wire wr_2559;
  wire wr_2560;
  wire wr_2561;
  wire wr_2562;
  wire wr_2563;
  wire wr_2564;
  wire wr_2565;
  wire wr_2566;
  wire wr_2567;
  wire wr_2568;
  wire wr_2569;
  wire wr_2570;
  wire wr_2571;
  wire wr_2572;
  wire wr_2573;
  wire wr_2574;
  wire wr_2575;
  wire wr_2576;
  wire wr_2577;
  wire wr_2578;
  wire wr_2579;
  wire wr_2580;
  wire wr_2581;
  wire wr_2582;
  wire wr_2583;
  wire wr_2584;
  wire wr_2585;
  wire wr_2586;
  wire wr_2587;
  wire wr_2588;
  wire wr_2589;
  wire wr_2590;
  wire wr_2591;
  wire wr_2592;
  wire wr_2593;
  wire wr_2594;
  wire wr_2595;
  wire wr_2596;
  wire wr_2597;
  wire wr_2598;
  wire wr_2599;
  wire wr_2600;
  wire wr_2601;
  wire wr_2602;
  wire wr_2603;
  wire wr_2604;
  wire wr_2605;
  wire wr_2606;
  wire wr_2607;
  wire wr_2608;
  wire wr_2609;
  wire wr_2610;
  wire wr_2611;
  wire wr_2612;
  wire wr_2613;
  wire wr_2614;
  wire wr_2615;
  wire wr_2616;
  wire wr_2617;
  wire wr_2618;
  wire wr_2619;
  wire wr_2620;
  wire wr_2621;
  wire wr_2622;
  wire wr_2623;
  wire wr_2624;
  wire wr_2625;
  wire wr_2626;
  wire wr_2627;
  wire wr_2628;
  wire wr_2629;
  wire wr_2630;
  wire wr_2631;
  wire wr_2632;
  wire wr_2633;
  wire wr_2634;
  wire wr_2635;
  wire wr_2636;
  wire wr_2637;
  wire wr_2638;
  wire wr_2639;
  wire wr_2640;
  wire wr_2641;
  wire wr_2642;
  wire wr_2643;
  wire wr_2644;
  wire wr_2645;
  wire wr_2646;
  wire wr_2647;
  wire wr_2648;
  wire wr_2649;
  wire wr_2650;
  wire wr_2651;
  wire wr_2652;
  wire wr_2653;
  wire wr_2654;
  wire wr_2655;
  wire wr_2656;
  wire wr_2657;
  wire wr_2658;
  wire wr_2659;
  wire wr_2660;
  wire wr_2661;
  wire wr_2662;
  wire wr_2663;
  wire wr_2664;
  wire wr_2665;
  wire wr_2666;
  wire wr_2667;
  wire wr_2668;
  wire wr_2669;
  wire wr_2670;
  wire wr_2671;
  wire wr_2672;
  wire wr_2673;
  wire wr_2674;
  wire wr_2675;
  wire wr_2676;
  wire wr_2677;
  wire wr_2678;
  wire wr_2679;
  wire wr_2680;
  wire wr_2681;
  wire wr_2682;
  wire wr_2683;
  wire wr_2684;
  wire wr_2685;
  wire wr_2686;
  wire wr_2687;
  wire wr_2688;
  wire wr_2689;
  wire wr_2690;
  wire wr_2691;
  wire wr_2692;
  wire wr_2693;
  wire wr_2694;
  wire wr_2695;
  wire wr_2696;
  wire wr_2697;
  wire wr_2698;
  wire wr_2699;
  wire wr_2700;
  wire wr_2701;
  wire wr_2702;
  wire wr_2703;
  wire wr_2704;
  wire wr_2705;
  wire wr_2706;
  wire wr_2707;
  wire wr_2708;
  wire wr_2709;
  wire wr_2710;
  wire wr_2711;
  wire wr_2712;
  wire wr_2713;
  wire wr_2714;
  wire wr_2715;
  wire wr_2716;
  wire wr_2717;
  wire wr_2718;
  wire wr_2719;
  wire wr_2720;
  wire wr_2721;
  wire wr_2722;
  wire wr_2723;
  wire wr_2724;
  wire wr_2725;
  wire wr_2726;
  wire wr_2727;
  wire wr_2728;
  wire wr_2729;
  wire wr_2730;
  wire wr_2731;
  wire wr_2732;
  wire wr_2733;
  wire wr_2734;
  wire wr_2735;
  wire wr_2736;
  wire wr_2737;
  wire wr_2738;
  wire wr_2739;
  wire wr_2740;
  wire wr_2741;
  wire wr_2742;
  wire wr_2743;
  wire wr_2744;
  wire wr_2745;
  wire wr_2746;
  wire wr_2747;
  wire wr_2748;
  wire wr_2749;
  wire wr_2750;
  wire wr_2751;
  wire wr_2752;
  wire wr_2753;
  wire wr_2754;
  wire wr_2755;
  wire wr_2756;
  wire wr_2757;
  wire wr_2758;
  wire wr_2759;
  wire wr_2760;
  wire wr_2761;
  wire wr_2762;
  wire wr_2763;
  wire wr_2764;
  wire wr_2765;
  wire wr_2766;
  wire wr_2767;
  wire wr_2768;
  wire wr_2769;
  wire wr_2770;
  wire wr_2771;
  wire wr_2772;
  wire wr_2773;
  wire wr_2774;
  wire wr_2775;
  wire wr_2776;
  wire wr_2777;
  wire wr_2778;
  wire wr_2779;
  wire wr_2780;
  wire wr_2781;
  wire wr_2782;
  wire wr_2783;
  wire wr_2784;
  wire wr_2785;
  wire wr_2786;
  wire wr_2787;
  wire wr_2788;
  wire wr_2789;
  wire wr_2790;
  wire wr_2791;
  wire wr_2792;
  wire wr_2793;
  wire wr_2794;
  wire wr_2795;
  wire wr_2796;
  wire wr_2797;
  wire wr_2798;
  wire wr_2799;
  wire wr_2800;
  wire wr_2801;
  wire wr_2802;
  wire wr_2803;
  wire wr_2804;
  wire wr_2805;
  wire wr_2806;
  wire wr_2807;
  wire wr_2808;
  wire wr_2809;
  wire wr_2810;
  wire wr_2811;
  wire wr_2812;
  wire wr_2813;
  wire wr_2814;
  wire wr_2815;
  wire wr_2816;
  wire wr_2817;
  wire wr_2818;
  wire wr_2819;
  wire wr_2820;
  wire wr_2821;
  wire wr_2822;
  wire wr_2823;
  wire wr_2824;
  wire wr_2825;
  wire wr_2826;
  wire wr_2827;
  wire wr_2828;
  wire wr_2829;
  wire wr_2830;
  wire wr_2831;
  wire wr_2832;
  wire wr_2833;
  wire wr_2834;
  wire wr_2835;
  wire wr_2836;
  wire wr_2837;
  wire wr_2838;
  wire wr_2839;
  wire wr_2840;
  wire wr_2841;
  wire wr_2842;
  wire wr_2843;
  wire wr_2844;
  wire wr_2845;
  wire wr_2846;
  wire wr_2847;
  wire wr_2848;
  wire wr_2849;
  wire wr_2850;
  wire wr_2851;
  wire wr_2852;
  wire wr_2853;
  wire wr_2854;
  wire wr_2855;
  wire wr_2856;
  wire wr_2857;
  wire wr_2858;
  wire wr_2859;
  wire wr_2860;
  wire wr_2861;
  wire wr_2862;
  wire wr_2863;
  wire wr_2864;
  wire wr_2865;
  wire wr_2866;
  wire wr_2867;
  wire wr_2868;
  wire wr_2869;
  wire wr_2870;
  wire wr_2871;
  wire wr_2872;
  wire wr_2873;
  wire wr_2874;
  wire wr_2875;
  wire wr_2876;
  wire wr_2877;
  wire wr_2878;
  wire wr_2879;
  wire wr_2880;
  wire wr_2881;
  wire wr_2882;
  wire wr_2883;
  wire wr_2884;
  wire wr_2885;
  wire wr_2886;
  wire wr_2887;
  wire wr_2888;
  wire wr_2889;
  wire wr_2890;
  wire wr_2891;
  wire wr_2892;
  wire wr_2893;
  wire wr_2894;
  wire wr_2895;
  wire wr_2896;
  wire wr_2897;
  wire wr_2898;
  wire wr_2899;
  wire wr_2900;
  wire wr_2901;
  wire wr_2902;
  wire wr_2903;
  wire wr_2904;
  wire wr_2905;
  wire wr_2906;
  wire wr_2907;
  wire wr_2908;
  wire wr_2909;
  wire wr_2910;
  wire wr_2911;
  wire wr_2912;
  wire wr_2913;
  wire wr_2914;
  wire wr_2915;
  wire wr_2916;
  wire wr_2917;
  wire wr_2918;
  wire wr_2919;
  wire wr_2920;
  wire wr_2921;
  wire wr_2922;
  wire wr_2923;
  wire wr_2924;
  wire wr_2925;
  wire wr_2926;
  wire wr_2927;
  wire wr_2928;
  wire wr_2929;
  wire wr_2930;
  wire wr_2931;
  wire wr_2932;
  wire wr_2933;
  wire wr_2934;
  wire wr_2935;
  wire wr_2936;
  wire wr_2937;
  wire wr_2938;
  wire wr_2939;
  wire wr_2940;
  wire wr_2941;
  wire wr_2942;
  wire wr_2943;
  wire wr_2944;
  wire wr_2945;
  wire wr_2946;
  wire wr_2947;
  wire wr_2948;
  wire wr_2949;
  wire wr_2950;
  wire wr_2951;
  wire wr_2952;
  wire wr_2953;
  wire wr_2954;
  wire wr_2955;
  wire wr_2956;
  wire wr_2957;
  wire wr_2958;
  wire wr_2959;
  wire wr_2960;
  wire wr_2961;
  wire wr_2962;
  wire wr_2963;
  wire wr_2964;
  wire wr_2965;
  wire wr_2966;
  wire wr_2967;
  wire wr_2968;
  wire wr_2969;
  wire wr_2970;
  wire wr_2971;
  wire wr_2972;
  wire wr_2973;
  wire wr_2974;
  wire wr_2975;
  wire wr_2976;
  wire wr_2977;
  wire wr_2978;
  wire wr_2979;
  wire wr_2980;
  wire wr_2981;
  wire wr_2982;
  wire wr_2983;
  wire wr_2984;
  wire wr_2985;
  wire wr_2986;
  wire wr_2987;
  wire wr_2988;
  wire wr_2989;
  wire wr_2990;
  wire wr_2991;
  wire wr_2992;
  wire wr_2993;
  wire wr_2994;
  wire wr_2995;
  wire wr_2996;
  wire wr_2997;
  wire wr_2998;
  wire wr_2999;
  wire wr_3000;
  wire wr_3001;
  wire wr_3002;
  wire wr_3003;
  wire wr_3004;
  wire wr_3005;
  wire wr_3006;
  wire wr_3007;
  wire wr_3008;
  wire wr_3009;
  wire wr_3010;
  wire wr_3011;
  wire wr_3012;
  wire wr_3013;
  wire wr_3014;
  wire wr_3015;
  wire wr_3016;
  wire wr_3017;
  wire wr_3018;
  wire wr_3019;
  wire wr_3020;
  wire wr_3021;
  wire wr_3022;
  wire wr_3023;
  wire wr_3024;
  wire wr_3025;
  wire wr_3026;
  wire wr_3027;
  wire wr_3028;
  wire wr_3029;
  wire wr_3030;
  wire wr_3031;
  wire wr_3032;
  wire wr_3033;
  wire wr_3034;
  wire wr_3035;
  wire wr_3036;
  wire wr_3037;
  wire wr_3038;
  wire wr_3039;
  wire wr_3040;
  wire wr_3041;
  wire wr_3042;
  wire wr_3043;
  wire wr_3044;
  wire wr_3045;
  wire wr_3046;
  wire wr_3047;
  wire wr_3048;
  wire wr_3049;
  wire wr_3050;
  wire wr_3051;
  wire wr_3052;
  wire wr_3053;
  wire wr_3054;
  wire wr_3055;
  wire wr_3056;
  wire wr_3057;
  wire wr_3058;
  wire wr_3059;
  wire wr_3060;
  wire wr_3061;
  wire wr_3062;
  wire wr_3063;
  wire wr_3064;
  wire wr_3065;
  wire wr_3066;
  wire wr_3067;
  wire wr_3068;
  wire wr_3069;
  wire wr_3070;
  wire wr_3071;
  wire wr_3072;
  wire wr_3073;
  wire wr_3074;
  wire wr_3075;
  wire wr_3076;
  wire wr_3077;
  wire wr_3078;
  wire wr_3079;
  wire wr_3080;
  wire wr_3081;
  wire wr_3082;
  wire wr_3083;
  wire wr_3084;
  wire wr_3085;
  wire wr_3086;
  wire wr_3087;
  wire wr_3088;
  wire wr_3089;
  wire wr_3090;
  wire wr_3091;
  wire wr_3092;
  wire wr_3093;
  wire wr_3094;
  wire wr_3095;
  wire wr_3096;
  wire wr_3097;
  wire wr_3098;
  wire wr_3099;
  wire wr_3100;
  wire wr_3101;
  wire wr_3102;
  wire wr_3103;
  wire wr_3104;
  wire wr_3105;
  wire wr_3106;
  wire wr_3107;
  wire wr_3108;
  wire wr_3109;
  wire wr_3110;
  wire wr_3111;
  wire wr_3112;
  wire wr_3113;
  wire wr_3114;
  wire wr_3115;
  wire wr_3116;
  wire wr_3117;
  wire wr_3118;
  wire wr_3119;
  wire wr_3120;
  wire wr_3121;
  wire wr_3122;
  wire wr_3123;
  wire wr_3124;
  wire wr_3125;
  wire wr_3126;
  wire wr_3127;
  wire wr_3128;
  wire wr_3129;
  wire wr_3130;
  wire wr_3131;
  wire wr_3132;
  wire wr_3133;
  wire wr_3134;
  wire wr_3135;
  wire wr_3136;
  wire wr_3137;
  wire wr_3138;
  wire wr_3139;
  wire wr_3140;
  wire wr_3141;
  wire wr_3142;
  wire wr_3143;
  wire wr_3144;
  wire wr_3145;
  wire wr_3146;
  wire wr_3147;
  wire wr_3148;
  wire wr_3149;
  wire wr_3150;
  wire wr_3151;
  wire wr_3152;
  wire wr_3153;
  wire wr_3154;
  wire wr_3155;
  wire wr_3156;
  wire wr_3157;
  wire wr_3158;
  wire wr_3159;
  wire wr_3160;
  wire wr_3161;
  wire wr_3162;
  wire wr_3163;
  wire wr_3164;
  wire wr_3165;
  wire wr_3166;
  wire wr_3167;
  wire wr_3168;
  wire wr_3169;
  wire wr_3170;
  wire wr_3171;
  wire wr_3172;
  wire wr_3173;
  wire wr_3174;
  wire wr_3175;
  wire wr_3176;
  wire wr_3177;
  wire wr_3178;
  wire wr_3179;
  wire wr_3180;
  wire wr_3181;
  wire wr_3182;
  wire wr_3183;
  wire wr_3184;
  wire wr_3185;
  wire wr_3186;
  wire wr_3187;
  wire wr_3188;
  wire wr_3189;
  wire wr_3190;
  wire wr_3191;
  wire wr_3192;
  wire wr_3193;
  wire wr_3194;
  wire wr_3195;
  wire wr_3196;
  wire wr_3197;
  wire wr_3198;
  wire wr_3199;
  wire wr_3200;
  wire wr_3201;
  wire wr_3202;
  wire wr_3203;
  wire wr_3204;
  wire wr_3205;
  wire wr_3206;
  wire wr_3207;
  wire wr_3208;
  wire wr_3209;
  wire wr_3210;
  wire wr_3211;
  wire wr_3212;
  wire wr_3213;
  wire wr_3214;
  wire wr_3215;
  wire wr_3216;
  wire wr_3217;
  wire wr_3218;
  wire wr_3219;
  wire wr_3220;
  wire wr_3221;
  wire wr_3222;
  wire wr_3223;
  wire wr_3224;
  wire wr_3225;
  wire wr_3226;
  wire wr_3227;
  wire wr_3228;
  wire wr_3229;
  wire wr_3230;
  wire wr_3231;
  wire wr_3232;
  wire wr_3233;
  wire wr_3234;
  wire wr_3235;
  wire wr_3236;
  wire wr_3237;
  wire wr_3238;
  wire wr_3239;
  wire wr_3240;
  wire wr_3241;
  wire wr_3242;
  wire wr_3243;
  wire wr_3244;
  wire wr_3245;
  wire wr_3246;
  wire wr_3247;
  wire wr_3248;
  wire wr_3249;
  wire wr_3250;
  wire wr_3251;
  wire wr_3252;
  wire wr_3253;
  wire wr_3254;
  wire wr_3255;
  wire wr_3256;
  wire wr_3257;
  wire wr_3258;
  wire wr_3259;
  wire wr_3260;
  wire wr_3261;
  wire wr_3262;
  wire wr_3263;
  wire wr_3264;
  wire wr_3265;
  wire wr_3266;
  wire wr_3267;
  wire wr_3268;
  wire wr_3269;
  wire wr_3270;
  wire wr_3271;
  wire wr_3272;
  wire wr_3273;
  wire wr_3274;
  wire wr_3275;
  wire wr_3276;
  wire wr_3277;
  wire wr_3278;
  wire wr_3279;
  wire wr_3280;
  wire wr_3281;
  wire wr_3282;
  wire wr_3283;
  wire wr_3284;
  wire wr_3285;
  wire wr_3286;
  wire wr_3287;
  wire wr_3288;
  wire wr_3289;
  wire wr_3290;
  wire wr_3291;
  wire wr_3292;
  wire wr_3293;
  wire wr_3294;
  wire wr_3295;
  wire wr_3296;
  wire wr_3297;
  wire wr_3298;
  wire wr_3299;
  wire wr_3300;
  wire wr_3301;
  wire wr_3302;
  wire wr_3303;
  wire wr_3304;
  wire wr_3305;
  wire wr_3306;
  wire wr_3307;
  wire wr_3308;
  wire wr_3309;
  wire wr_3310;
  wire wr_3311;
  wire wr_3312;
  wire wr_3313;
  wire wr_3314;
  wire wr_3315;
  wire wr_3316;
  wire wr_3317;
  wire wr_3318;
  wire wr_3319;
  wire wr_3320;
  wire wr_3321;
  wire wr_3322;
  wire wr_3323;
  wire wr_3324;
  wire wr_3325;
  wire wr_3326;
  wire wr_3327;
  wire wr_3328;
  wire wr_3329;
  wire wr_3330;
  wire wr_3331;
  wire wr_3332;
  wire wr_3333;
  wire wr_3334;
  wire wr_3335;
  wire wr_3336;
  wire wr_3337;
  wire wr_3338;
  wire wr_3339;
  wire wr_3340;
  wire wr_3341;
  wire wr_3342;
  wire wr_3343;
  wire wr_3344;
  wire wr_3345;
  wire wr_3346;
  wire wr_3347;
  wire wr_3348;
  wire wr_3349;
  wire wr_3350;
  wire wr_3351;
  wire wr_3352;
  wire wr_3353;
  wire wr_3354;
  wire wr_3355;
  wire wr_3356;
  wire wr_3357;
  wire wr_3358;
  wire wr_3359;
  wire wr_3360;
  wire wr_3361;
  wire wr_3362;
  wire wr_3363;
  wire wr_3364;
  wire wr_3365;
  wire wr_3366;
  wire wr_3367;
  wire wr_3368;
  wire wr_3369;
  wire wr_3370;
  wire wr_3371;
  wire wr_3372;
  wire wr_3373;
  wire wr_3374;
  wire wr_3375;
  wire wr_3376;
  wire wr_3377;
  wire wr_3378;
  wire wr_3379;
  wire wr_3380;
  wire wr_3381;
  wire wr_3382;
  wire wr_3383;
  wire wr_3384;
  wire wr_3385;
  wire wr_3386;
  wire wr_3387;
  wire wr_3388;
  wire wr_3389;
  wire wr_3390;
  wire wr_3391;
  wire wr_3392;
  wire wr_3393;
  wire wr_3394;
  wire wr_3395;

  not    g1( wr_154  ,           G41     );
  not    g2( wr_157  ,           G3701   );
  not    g3( wr_184  ,           G1462   );
  not    g4( wr_185  ,           G9      );
  not    g5( wr_186  ,           G12     );
  not    g6( wr_188  ,           G18     );
  not    g7( wr_195  ,           G1480   );
  not    g8( wr_202  ,           G106    );
  not    g9( wr_209  ,           G1469   );
  not   g10( wr_247  ,           G2247   );
  not   g11( wr_254  ,           G2253   );
  not   g12( wr_279  ,           G2239   );
  not   g13( wr_289  ,           G2236   );
  not   g14( wr_296  ,           G135    );
  not   g15( wr_298  ,           G158    );
  not   g16( wr_305  ,           G2230   );
  not   g17( wr_310  ,           G144    );
  not   g18( wr_312  ,           G159    );
  not   g19( wr_320  ,           G2224   );
  not   g20( wr_325  ,           G2218   );
  not   g21( wr_326  ,           G138    );
  not   g22( wr_328  ,           G160    );
  not   g23( wr_335  ,           G147    );
  not   g24( wr_337  ,           G151    );
  not   g25( wr_407  ,           G2211   );
  not   g26( wr_423  ,           G219    );
  not   g27( wr_425  ,           G66     );
  not   g28( wr_432  ,           G220    );
  not   g29( wr_434  ,           G50     );
  not   g30( wr_441  ,           G4427   );
  not   g31( wr_442  ,           G221    );
  not   g32( wr_444  ,           G32     );
  not   g33( wr_451  ,           G4432   );
  not   g34( wr_456  ,           G222    );
  not   g35( wr_458  ,           G35     );
  not   g36( wr_479  ,           G4420   );
  not   g37( wr_490  ,           G4415   );
  not   g38( wr_491  ,           G223    );
  not   g39( wr_493  ,           G47     );
  not   g40( wr_500  ,           G224    );
  not   g41( wr_502  ,           G121    );
  not   g42( wr_509  ,           G4410   );
  not   g43( wr_514  ,           G225    );
  not   g44( wr_516  ,           G94     );
  not   g45( wr_524  ,           G4405   );
  not   g46( wr_529  ,           G4400   );
  not   g47( wr_530  ,           G226    );
  not   g48( wr_532  ,           G97     );
  not   g49( wr_539  ,           G217    );
  not   g50( wr_541  ,           G118    );
  not   g51( wr_572  ,           G3729   );
  not   g52( wr_573  ,           G234    );
  not   g53( wr_575  ,           G130    );
  not   g54( wr_582  ,           G3743   );
  not   g55( wr_583  ,           G232    );
  not   g56( wr_585  ,           G124    );
  not   g57( wr_602  ,           G3737   );
  not   g58( wr_603  ,           G233    );
  not   g59( wr_605  ,           G127    );
  not   g60( wr_618  ,           G3717   );
  not   g61( wr_619  ,           G236    );
  not   g62( wr_621  ,           G23     );
  not   g63( wr_628  ,           G3711   );
  not   g64( wr_629  ,           G237    );
  not   g65( wr_631  ,           G26     );
  not   g66( wr_638  ,           G3705   );
  not   g67( wr_639  ,           G238    );
  not   g68( wr_641  ,           G29     );
  not   g69( wr_648  ,           G3723   );
  not   g70( wr_649  ,           G235    );
  not   g71( wr_651  ,           G103    );
  not   g72( wr_668  ,           G4394   );
  not   g73( wr_593  ,           G231    );
  not   g74( wr_595  ,           G100    );
  not   g75( wr_1313 ,           G205    );
  not   g76( wr_1317 ,           G75     );
  not   g77( wr_233  ,           G2256   );
  not   g78( wr_422  ,           G4437   );
  not   g79( wr_1301 ,           G204    );
  not   g80( wr_1305 ,           G73     );
  not   g81( wr_592  ,           G3749   );
  not   g82( wr_1270 ,           G207    );
  not   g83( wr_1274 ,           G74     );
  nor   g84( wr_1284 , G70     , G18     );
  not   g85( wr_906  ,           G64     );
  not   g86( wr_914  ,           G178    );
  not   g87( wr_917  ,           G85     );
  not   g88( wr_1124 ,           G193    );
  not   g89( wr_1128 ,           G80     );
  not   g90( wr_1136 ,           G194    );
  not   g91( wr_1140 ,           G81     );
  not   g92( wr_1252 ,           G201    );
  not   g93( wr_1256 ,           G55     );
  not   g94( wr_1289 ,           G206    );
  not   g95( wr_1293 ,           G76     );
  not   g96( wr_802  ,           G88     );
  not   g97( wr_813  ,           G112    );
  not   g98( wr_959  ,           G171    );
  not   g99( wr_962  ,           G65     );
  not  g100( wr_1228 ,           G203    );
  not  g101( wr_1232 ,           G53     );
  not  g102( wr_834  ,           G110    );
  not  g103( wr_845  ,           G109    );
  not  g104( wr_930  ,           G179    );
  not  g105( wr_933  ,           G84     );
  not  g106( wr_1048 ,           G189    );
  not  g107( wr_1052 ,           G62     );
  not  g108( wr_1060 ,           G190    );
  not  g109( wr_1064 ,           G61     );
  not  g110( wr_1152 ,           G195    );
  not  g111( wr_1156 ,           G59     );
  not  g112( wr_1169 ,           G196    );
  not  g113( wr_1181 ,           G187    );
  not  g114( wr_1185 ,           G77     );
  not  g115( wr_1216 ,           G202    );
  not  g116( wr_1220 ,           G54     );
  not  g117( wr_1750 ,           G229    );
  not  g118( wr_1755 ,           G239    );
  not  g119( wr_1757 ,           G44     );
  not  g120( wr_1806 ,           G227    );
  not  g121( wr_1808 ,           G115    );
  not  g122( wr_2166 ,           G198    );
  not  g123( wr_2170 ,           G208    );
  not  g124( wr_2219 ,           G197    );
  not  g125( wr_791  ,           G87     );
  not  g126( wr_947  ,           G180    );
  not  g127( wr_950  ,           G83     );
  not  g128( wr_216  ,           G1486   );
  not  g129( wr_871  ,           G63     );
  not  g130( wr_1088 ,           G192    );
  not  g131( wr_1092 ,           G79     );
  not  g132( wr_1173 ,           G78     );
  not  g133( wr_1240 ,           G200    );
  not  g134( wr_1244 ,           G56     );
  not  g135( wr_1965 ,           G69     );
  not  g136( wr_1968 ,           G70     );
  not  g137( wr_2020 ,           G58     );
  not  g138( wr_779  ,           G113    );
  not  g139( wr_771  ,           G111    );
  not  g140( wr_856  ,           G86     );
  not  g141( wr_1071 ,           G191    );
  not  g142( wr_1075 ,           G60     );
  not  g143( wr_1657 ,           G141    );
  not  g144( wr_1659 ,           G161    );
  not  g145( wr_1914 ,           G114    );
  not  g146( wr_2074 ,           G181    );
  not  g147( wr_169  ,           G1492   );
  not  g148( wr_170  ,           G4528   );
  not  g149( wr_176  ,           G1496   );
  not  g150( wr_1862 ,           G82     );
  not  g151( wr_164  ,           G4526   );
  not  g152( wr_168  ,           G38     );
  not  g153( wr_1893 ,           G1455   );
  not  g154( wr_1897 ,           G2204   );
  not  g155( wr_1335 ,           G89     );
  not  g156( wr_111  ,           G228    );
  not  g157( wr_112  ,           G240    );
  not  g158( wr_120  ,           G218    );
  not  g159( wr_121  ,           G230    );
  not  g160( wr_110  ,           G150    );
  not  g161( wr_119  ,           G210    );
  not  g162( wr_129  ,           G185    );
  not  g163( wr_130  ,           G186    );
  not  g164( wr_138  ,           G188    );
  not  g165( wr_139  ,           G199    );
  not  g166( wr_109  ,           G184    );
  not  g167( wr_118  ,           G152    );
  not  g168( wr_128  ,           G183    );
  not  g169( wr_137  ,           G162    );
  not  g170( wr_127  ,           G182    );
  not  g171( wr_136  ,           G172    );
  not  g172( wr_147  ,           G133    );
  not  g173( wr_148  ,           G134    );
  not  g174( wr_145  ,           G1197   );
  nor  g175( wr_108  , G57     , G5      );
  not  g176( wr_152  ,           G1      );
  not  g177( wr_153  ,           G163    );
  not  g178( G279    ,           G15     );
  not  g179( G2      ,           G1      );
  not  g180( G3      ,           G1      );
  not  g181( G450    ,           G1459   );
  not  g182( G448    ,           G1469   );
  not  g183( G444    ,           G1480   );
  not  g184( G442    ,           G1486   );
  not  g185( G440    ,           G1492   );
  not  g186( G438    ,           G1496   );
  not  g187( G496    ,           G2208   );
  not  g188( G494    ,           G2218   );
  not  g189( G492    ,           G2224   );
  not  g190( G490    ,           G2230   );
  not  g191( G488    ,           G2236   );
  not  g192( G486    ,           G2239   );
  not  g193( G484    ,           G2247   );
  not  g194( G482    ,           G2253   );
  not  g195( G480    ,           G2256   );
  not  g196( G560    ,           G3698   );
  not  g197( G542    ,           G3701   );
  not  g198( G558    ,           G3705   );
  not  g199( G556    ,           G3711   );
  not  g200( G554    ,           G3717   );
  not  g201( G552    ,           G3723   );
  not  g202( G550    ,           G3729   );
  not  g203( G548    ,           G3737   );
  not  g204( G546    ,           G3743   );
  not  g205( G544    ,           G3749   );
  not  g206( G540    ,           G4393   );
  not  g207( G538    ,           G4400   );
  not  g208( G536    ,           G4405   );
  not  g209( G534    ,           G4410   );
  not  g210( G532    ,           G4415   );
  not  g211( G530    ,           G4420   );
  not  g212( G528    ,           G4427   );
  not  g213( G526    ,           G4432   );
  not  g214( G524    ,           G4437   );
  not  g215( G436    ,           G1462   );
  not  g216( G478    ,           G2211   );
  not  g217( G522    ,           G4394   );
  not  g218( G432    ,           G1      );
  not  g219( G446    ,           G106    );
  not  g220( G286    ,           G15     );
  not  g221( G341    ,           G15     );
  not  g222( G453    ,           G1      );
  nor  g223( wr_155  , wr_154  , G18     );
  nor  g224( wr_158  , wr_157  , G18     );
  nor  g225( wr_187  , wr_186  , wr_185  );
  nor  g226( wr_189  , G209    , wr_188  );
  nor  g227( wr_196  , G214    , wr_188  );
  nor  g228( wr_203  , G215    , wr_188  );
  nor  g229( wr_210  , G216    , wr_188  );
  nor  g230( wr_234  , G153    , wr_188  );
  nor  g231( wr_240  , G154    , wr_188  );
  nor  g232( wr_248  , G155    , wr_188  );
  nor  g233( wr_258  , G156    , wr_188  );
  nor  g234( wr_290  , G157    , wr_188  );
  nor  g235( wr_297  , wr_296  , G18     );
  nor  g236( wr_299  , wr_298  , wr_188  );
  nor  g237( wr_311  , wr_310  , G18     );
  nor  g238( wr_313  , wr_312  , wr_188  );
  nor  g239( wr_327  , wr_326  , G18     );
  nor  g240( wr_329  , wr_328  , wr_188  );
  nor  g241( wr_336  , wr_335  , G18     );
  nor  g242( wr_338  , wr_337  , wr_188  );
  nor  g243( wr_424  , wr_423  , wr_188  );
  nor  g244( wr_426  , wr_425  , G18     );
  nor  g245( wr_433  , wr_432  , wr_188  );
  nor  g246( wr_435  , wr_434  , G18     );
  nor  g247( wr_443  , wr_442  , wr_188  );
  nor  g248( wr_445  , wr_444  , G18     );
  nor  g249( wr_457  , wr_456  , wr_188  );
  nor  g250( wr_459  , wr_458  , G18     );
  nor  g251( wr_492  , wr_491  , wr_188  );
  nor  g252( wr_494  , wr_493  , G18     );
  nor  g253( wr_501  , wr_500  , wr_188  );
  nor  g254( wr_503  , wr_502  , G18     );
  nor  g255( wr_515  , wr_514  , wr_188  );
  nor  g256( wr_517  , wr_516  , G18     );
  nor  g257( wr_531  , wr_530  , wr_188  );
  nor  g258( wr_533  , wr_532  , G18     );
  nor  g259( wr_540  , wr_539  , wr_188  );
  nor  g260( wr_542  , wr_541  , G18     );
  nor  g261( wr_574  , wr_573  , wr_188  );
  nor  g262( wr_576  , wr_575  , G18     );
  nor  g263( wr_584  , wr_583  , wr_188  );
  nor  g264( wr_586  , wr_585  , G18     );
  nor  g265( wr_604  , wr_603  , wr_188  );
  nor  g266( wr_606  , wr_605  , G18     );
  nor  g267( wr_620  , wr_619  , wr_188  );
  nor  g268( wr_622  , wr_621  , G18     );
  nor  g269( wr_630  , wr_629  , wr_188  );
  nor  g270( wr_632  , wr_631  , G18     );
  nor  g271( wr_640  , wr_639  , wr_188  );
  nor  g272( wr_642  , wr_641  , G18     );
  nor  g273( wr_650  , wr_649  , wr_188  );
  nor  g274( wr_652  , wr_651  , G18     );
  nor  g275( wr_594  , wr_593  , wr_188  );
  nor  g276( wr_596  , wr_595  , G18     );
  nor  g277( wr_1314 , wr_1313 , wr_188  );
  nor  g278( wr_1316 , G3717   , wr_188  );
  nor  g279( wr_1318 , wr_1317 , G18     );
  nor  g280( wr_1282 , wr_154  , G18     );
  nor  g281( wr_1302 , wr_1301 , wr_188  );
  nor  g282( wr_1304 , G3723   , wr_188  );
  nor  g283( wr_1306 , wr_1305 , G18     );
  nor  g284( wr_1271 , wr_1270 , wr_188  );
  nor  g285( wr_1273 , G3705   , wr_188  );
  nor  g286( wr_1275 , wr_1274 , G18     );
  nor  g287( wr_903  , G177    , wr_188  );
  nor  g288( wr_907  , wr_906  , G18     );
  nor  g289( wr_908  , G2236   , wr_188  );
  nor  g290( wr_915  , wr_914  , wr_188  );
  nor  g291( wr_918  , wr_917  , G18     );
  nor  g292( wr_919  , G2230   , wr_188  );
  nor  g293( wr_1125 , wr_1124 , wr_188  );
  nor  g294( wr_1127 , G4415   , wr_188  );
  nor  g295( wr_1129 , wr_1128 , G18     );
  nor  g296( wr_1137 , wr_1136 , wr_188  );
  nor  g297( wr_1139 , G4410   , wr_188  );
  nor  g298( wr_1141 , wr_1140 , G18     );
  nor  g299( wr_1253 , wr_1252 , wr_188  );
  nor  g300( wr_1255 , G3743   , wr_188  );
  nor  g301( wr_1257 , wr_1256 , G18     );
  nor  g302( wr_1290 , wr_1289 , wr_188  );
  nor  g303( wr_1292 , G3711   , wr_188  );
  nor  g304( wr_1294 , wr_1293 , G18     );
  nor  g305( wr_217  , G213    , wr_188  );
  nor  g306( wr_799  , G166    , wr_188  );
  nor  g307( wr_803  , wr_802  , G18     );
  nor  g308( wr_804  , G1486   , wr_188  );
  nor  g309( wr_810  , G167    , wr_188  );
  nor  g310( wr_814  , wr_813  , G18     );
  nor  g311( wr_815  , G1480   , wr_188  );
  nor  g312( wr_960  , wr_959  , wr_188  );
  nor  g313( wr_963  , wr_962  , G18     );
  nor  g314( wr_964  , G2211   , wr_188  );
  nor  g315( wr_1229 , wr_1228 , wr_188  );
  nor  g316( wr_1231 , G3729   , wr_188  );
  nor  g317( wr_1233 , wr_1232 , G18     );
  nor  g318( wr_831  , G173    , wr_188  );
  nor  g319( wr_835  , wr_834  , G18     );
  nor  g320( wr_836  , G2256   , wr_188  );
  nor  g321( wr_842  , G174    , wr_188  );
  nor  g322( wr_846  , wr_845  , G18     );
  nor  g323( wr_847  , G2253   , wr_188  );
  nor  g324( wr_931  , wr_930  , wr_188  );
  nor  g325( wr_934  , wr_933  , G18     );
  nor  g326( wr_935  , G2224   , wr_188  );
  nor  g327( wr_1049 , wr_1048 , wr_188  );
  nor  g328( wr_1051 , G4437   , wr_188  );
  nor  g329( wr_1053 , wr_1052 , G18     );
  nor  g330( wr_1061 , wr_1060 , wr_188  );
  nor  g331( wr_1063 , G4432   , wr_188  );
  nor  g332( wr_1065 , wr_1064 , G18     );
  nor  g333( wr_1153 , wr_1152 , wr_188  );
  nor  g334( wr_1155 , G4405   , wr_188  );
  nor  g335( wr_1157 , wr_1156 , G18     );
  nor  g336( wr_1170 , wr_1169 , wr_188  );
  nor  g337( wr_1182 , wr_1181 , wr_188  );
  nor  g338( wr_1184 , G4394   , wr_188  );
  nor  g339( wr_1186 , wr_1185 , G18     );
  nor  g340( wr_1217 , wr_1216 , wr_188  );
  nor  g341( wr_1219 , G3737   , wr_188  );
  nor  g342( wr_1221 , wr_1220 , G18     );
  nor  g343( wr_1751 , wr_1750 , wr_188  );
  nor  g344( wr_1752 , wr_154  , G18     );
  nor  g345( wr_1756 , wr_1755 , wr_188  );
  nor  g346( wr_1758 , wr_1757 , G18     );
  nor  g347( wr_1807 , wr_1806 , wr_188  );
  nor  g348( wr_1809 , wr_1808 , G18     );
  nor  g349( wr_2167 , wr_2166 , wr_188  );
  nor  g350( wr_2171 , wr_2170 , wr_188  );
  nor  g351( wr_2220 , wr_2219 , wr_188  );
  nor  g352( wr_788  , G168    , wr_188  );
  nor  g353( wr_792  , wr_791  , G18     );
  nor  g354( wr_793  , G106    , wr_188  );
  nor  g355( wr_948  , wr_947  , wr_188  );
  nor  g356( wr_951  , wr_950  , G18     );
  nor  g357( wr_952  , G2218   , wr_188  );
  nor  g358( wr_768  , G169    , wr_188  );
  nor  g359( wr_868  , G176    , wr_188  );
  nor  g360( wr_872  , wr_871  , G18     );
  nor  g361( wr_873  , G2239   , wr_188  );
  nor  g362( wr_1089 , wr_1088 , wr_188  );
  nor  g363( wr_1091 , G4420   , wr_188  );
  nor  g364( wr_1093 , wr_1092 , G18     );
  nor  g365( wr_1172 , G4400   , wr_188  );
  nor  g366( wr_1174 , wr_1173 , G18     );
  nor  g367( wr_1241 , wr_1240 , wr_188  );
  nor  g368( wr_1243 , G3749   , wr_188  );
  nor  g369( wr_1245 , wr_1244 , G18     );
  nor  g370( wr_1964 , G3698   , wr_188  );
  nor  g371( wr_1966 , wr_1965 , G18     );
  nor  g372( wr_1969 , wr_1968 , G18     );
  nor  g373( wr_1970 , G3701   , wr_188  );
  nor  g374( wr_2019 , G4393   , wr_188  );
  nor  g375( wr_2021 , wr_2020 , G18     );
  nor  g376( wr_780  , wr_779  , G18     );
  nor  g377( wr_781  , G1462   , wr_188  );
  nor  g378( wr_772  , wr_771  , G18     );
  nor  g379( wr_773  , G1469   , wr_188  );
  nor  g380( wr_853  , G175    , wr_188  );
  nor  g381( wr_857  , wr_856  , G18     );
  nor  g382( wr_858  , G2247   , wr_188  );
  nor  g383( wr_1072 , wr_1071 , wr_188  );
  nor  g384( wr_1074 , G4427   , wr_188  );
  nor  g385( wr_1076 , wr_1075 , G18     );
  nor  g386( wr_1658 , wr_1657 , G18     );
  nor  g387( wr_1660 , wr_1659 , wr_188  );
  nor  g388( wr_1915 , wr_1914 , G18     );
  nor  g389( wr_1916 , G1459   , wr_188  );
  nor  g390( wr_2075 , wr_2074 , wr_188  );
  nor  g391( wr_2121 , G170    , wr_188  );
  nor  g392( wr_171  , wr_170  , wr_169  );
  nor  g393( wr_177  , wr_170  , wr_176  );
  nor  g394( wr_756  , wr_170  , G1455   );
  nor  g395( wr_761  , wr_170  , G2204   );
  nor  g396( wr_1863 , wr_1862 , G18     );
  nor  g397( wr_1864 , G2208   , wr_188  );
  not  g398( wr_1285 ,           wr_1284 );
  nor  g399( wr_1689 , G212    , wr_188  );
  nor  g400( wr_1692 , G211    , wr_188  );
  nor  g401( wr_2104 , G165    , wr_188  );
  nor  g402( wr_2107 , G164    , wr_188  );
  nor  g403( wr_1894 , wr_1893 , G18     );
  nor  g404( wr_1895 , G1492   , wr_188  );
  nor  g405( wr_1898 , wr_1897 , G18     );
  nor  g406( wr_1899 , G1496   , wr_188  );
  nor  g407( wr_113  , wr_112  , wr_111  );
  nor  g408( wr_122  , wr_121  , wr_120  );
  nor  g409( wr_131  , wr_130  , wr_129  );
  nor  g410( wr_140  , wr_139  , wr_138  );
  nor  g411( wr_149  , wr_148  , wr_147  );
  nor  g412( wr_146  , wr_145  , G5      );
  not  g413( G402    ,           wr_108  );
  nor  g414( G278    , wr_153  , wr_152  );
  not  g415( wr_156  ,           wr_155  );
  not  g416( wr_159  ,           wr_158  );
  nor  g417( wr_161  , wr_158  , wr_155  );
  nor  g418( wr_190  , wr_189  , wr_187  );
  nor  g419( wr_197  , wr_196  , wr_187  );
  nor  g420( wr_204  , wr_203  , wr_187  );
  nor  g421( wr_211  , wr_210  , wr_187  );
  nor  g422( wr_241  , wr_240  , wr_187  );
  nor  g423( wr_249  , wr_248  , wr_187  );
  nor  g424( wr_259  , wr_258  , wr_187  );
  nor  g425( wr_291  , wr_290  , wr_187  );
  nor  g426( wr_300  , wr_299  , wr_297  );
  nor  g427( wr_314  , wr_313  , wr_311  );
  nor  g428( wr_330  , wr_329  , wr_327  );
  nor  g429( wr_339  , wr_338  , wr_336  );
  nor  g430( wr_436  , wr_435  , wr_433  );
  nor  g431( wr_446  , wr_445  , wr_443  );
  nor  g432( wr_460  , wr_459  , wr_457  );
  nor  g433( wr_495  , wr_494  , wr_492  );
  nor  g434( wr_504  , wr_503  , wr_501  );
  nor  g435( wr_518  , wr_517  , wr_515  );
  nor  g436( wr_534  , wr_533  , wr_531  );
  nor  g437( wr_543  , wr_542  , wr_540  );
  nor  g438( wr_577  , wr_576  , wr_574  );
  nor  g439( wr_587  , wr_586  , wr_584  );
  nor  g440( wr_607  , wr_606  , wr_604  );
  nor  g441( wr_623  , wr_622  , wr_620  );
  nor  g442( wr_633  , wr_632  , wr_630  );
  nor  g443( wr_643  , wr_642  , wr_640  );
  nor  g444( wr_653  , wr_652  , wr_650  );
  nor  g445( wr_235  , wr_234  , wr_187  );
  nor  g446( wr_427  , wr_426  , wr_424  );
  nor  g447( wr_597  , wr_596  , wr_594  );
  nor  g448( wr_1315 , wr_1314 , wr_622  );
  nor  g449( wr_1319 , wr_1318 , wr_1316 );
  not  g450( wr_1283 ,           wr_1282 );
  nor  g451( wr_1303 , wr_1302 , wr_652  );
  nor  g452( wr_1307 , wr_1306 , wr_1304 );
  nor  g453( wr_1272 , wr_1271 , wr_642  );
  nor  g454( wr_1276 , wr_1275 , wr_1273 );
  nor  g455( wr_904  , wr_903  , wr_187  );
  nor  g456( wr_909  , wr_908  , wr_907  );
  nor  g457( wr_916  , wr_915  , wr_297  );
  nor  g458( wr_920  , wr_919  , wr_918  );
  nor  g459( wr_1126 , wr_1125 , wr_494  );
  nor  g460( wr_1130 , wr_1129 , wr_1127 );
  nor  g461( wr_1138 , wr_1137 , wr_503  );
  nor  g462( wr_1142 , wr_1141 , wr_1139 );
  nor  g463( wr_1254 , wr_1253 , wr_586  );
  nor  g464( wr_1258 , wr_1257 , wr_1255 );
  nor  g465( wr_1291 , wr_1290 , wr_632  );
  nor  g466( wr_1295 , wr_1294 , wr_1292 );
  nor  g467( wr_218  , wr_217  , wr_187  );
  nor  g468( wr_800  , wr_799  , wr_187  );
  nor  g469( wr_805  , wr_804  , wr_803  );
  nor  g470( wr_811  , wr_810  , wr_187  );
  nor  g471( wr_816  , wr_815  , wr_814  );
  nor  g472( wr_961  , wr_960  , wr_336  );
  nor  g473( wr_965  , wr_964  , wr_963  );
  nor  g474( wr_1230 , wr_1229 , wr_576  );
  nor  g475( wr_1234 , wr_1233 , wr_1231 );
  nor  g476( wr_832  , wr_831  , wr_187  );
  nor  g477( wr_837  , wr_836  , wr_835  );
  nor  g478( wr_843  , wr_842  , wr_187  );
  nor  g479( wr_848  , wr_847  , wr_846  );
  nor  g480( wr_932  , wr_931  , wr_311  );
  nor  g481( wr_936  , wr_935  , wr_934  );
  nor  g482( wr_1050 , wr_1049 , wr_426  );
  nor  g483( wr_1054 , wr_1053 , wr_1051 );
  nor  g484( wr_1062 , wr_1061 , wr_435  );
  nor  g485( wr_1066 , wr_1065 , wr_1063 );
  nor  g486( wr_1154 , wr_1153 , wr_517  );
  nor  g487( wr_1158 , wr_1157 , wr_1155 );
  nor  g488( wr_1171 , wr_1170 , wr_533  );
  nor  g489( wr_1183 , wr_1182 , wr_542  );
  nor  g490( wr_1187 , wr_1186 , wr_1184 );
  nor  g491( wr_1218 , wr_1217 , wr_606  );
  nor  g492( wr_1222 , wr_1221 , wr_1219 );
  nor  g493( wr_1753 , wr_1752 , wr_1751 );
  nor  g494( wr_1759 , wr_1758 , wr_1756 );
  nor  g495( wr_1810 , wr_1809 , wr_1807 );
  nor  g496( wr_2168 , wr_2167 , wr_1752 );
  nor  g497( wr_2172 , wr_2171 , wr_1758 );
  nor  g498( wr_2221 , wr_2220 , wr_1809 );
  nor  g499( wr_789  , wr_788  , wr_187  );
  nor  g500( wr_794  , wr_793  , wr_792  );
  nor  g501( wr_949  , wr_948  , wr_327  );
  nor  g502( wr_953  , wr_952  , wr_951  );
  nor  g503( wr_769  , wr_768  , wr_187  );
  nor  g504( wr_869  , wr_868  , wr_187  );
  nor  g505( wr_874  , wr_873  , wr_872  );
  nor  g506( wr_1090 , wr_1089 , wr_459  );
  nor  g507( wr_1094 , wr_1093 , wr_1091 );
  nor  g508( wr_1175 , wr_1174 , wr_1172 );
  nor  g509( wr_1242 , wr_1241 , wr_596  );
  nor  g510( wr_1246 , wr_1245 , wr_1243 );
  nor  g511( wr_1967 , wr_1966 , wr_1964 );
  nor  g512( wr_1971 , wr_1970 , wr_1969 );
  nor  g513( wr_2022 , wr_2021 , wr_2019 );
  nor  g514( wr_782  , wr_781  , wr_780  );
  nor  g515( wr_774  , wr_773  , wr_772  );
  not  g516( wr_785  ,           wr_187  );
  nor  g517( wr_854  , wr_853  , wr_187  );
  nor  g518( wr_859  , wr_858  , wr_857  );
  nor  g519( wr_1073 , wr_1072 , wr_445  );
  nor  g520( wr_1077 , wr_1076 , wr_1074 );
  nor  g521( wr_1661 , wr_1660 , wr_1658 );
  not  g522( wr_1706 ,           wr_189  );
  nor  g523( wr_1917 , wr_1916 , wr_1915 );
  nor  g524( wr_2076 , wr_2075 , wr_1658 );
  not  g525( wr_2122 ,           wr_2121 );
  not  g526( wr_172  ,           wr_171  );
  not  g527( wr_178  ,           wr_177  );
  not  g528( wr_757  ,           wr_756  );
  not  g529( wr_762  ,           wr_761  );
  nor  g530( wr_1865 , wr_1864 , wr_1863 );
  nor  g531( wr_174  , wr_171  , G38     );
  nor  g532( wr_180  , wr_177  , G38     );
  nor  g533( wr_759  , wr_756  , G38     );
  nor  g534( wr_764  , wr_761  , G38     );
  nor  g535( wr_1287 , wr_1284 , wr_1282 );
  nor  g536( wr_1690 , wr_1689 , wr_187  );
  nor  g537( wr_1693 , wr_1692 , wr_187  );
  nor  g538( wr_2105 , wr_2104 , wr_187  );
  nor  g539( wr_2108 , wr_2107 , wr_187  );
  nor  g540( wr_1896 , wr_1895 , wr_1894 );
  nor  g541( wr_1900 , wr_1899 , wr_1898 );
  nor  g542( wr_3001 , wr_171  , wr_168  );
  not  g543( wr_114  ,           wr_113  );
  not  g544( wr_123  ,           wr_122  );
  nor  g545( wr_367  , wr_171  , wr_168  );
  nor  g546( wr_993  , wr_756  , wr_168  );
  not  g547( wr_132  ,           wr_131  );
  not  g548( wr_141  ,           wr_140  );
  nor  g549( wr_366  , wr_177  , wr_168  );
  nor  g550( wr_992  , wr_761  , wr_168  );
  not  g551( wr_150  ,           wr_149  );
  not  g552( G284    ,           wr_146  );
  not  g553( G289    ,           wr_146  );
  nor  g554( wr_160  , wr_159  , wr_156  );
  not  g555( wr_191  ,           wr_190  );
  nor  g556( wr_193  , wr_190  , G1462   );
  not  g557( wr_198  ,           wr_197  );
  nor  g558( wr_200  , wr_197  , G1480   );
  not  g559( wr_205  ,           wr_204  );
  nor  g560( wr_207  , wr_204  , G106    );
  not  g561( wr_212  ,           wr_211  );
  nor  g562( wr_214  , wr_211  , G1469   );
  not  g563( wr_242  ,           wr_241  );
  not  g564( wr_250  ,           wr_249  );
  not  g565( wr_260  ,           wr_259  );
  not  g566( wr_292  ,           wr_291  );
  nor  g567( wr_306  , wr_300  , wr_305  );
  not  g568( wr_307  ,           wr_300  );
  nor  g569( wr_321  , wr_314  , wr_320  );
  not  g570( wr_322  ,           wr_314  );
  nor  g571( wr_331  , wr_330  , wr_325  );
  not  g572( wr_332  ,           wr_330  );
  nor  g573( wr_340  , wr_339  , G2211   );
  nor  g574( wr_408  , wr_339  , wr_407  );
  not  g575( wr_409  ,           wr_339  );
  not  g576( wr_448  ,           wr_446  );
  not  g577( wr_453  ,           wr_436  );
  not  g578( wr_481  ,           wr_460  );
  not  g579( wr_497  ,           wr_495  );
  nor  g580( wr_510  , wr_504  , wr_509  );
  not  g581( wr_511  ,           wr_504  );
  nor  g582( wr_525  , wr_518  , wr_524  );
  not  g583( wr_526  ,           wr_518  );
  nor  g584( wr_535  , wr_534  , wr_529  );
  not  g585( wr_536  ,           wr_534  );
  nor  g586( wr_544  , wr_543  , G4394   );
  not  g587( wr_579  ,           wr_577  );
  not  g588( wr_589  ,           wr_587  );
  not  g589( wr_609  ,           wr_607  );
  nor  g590( wr_624  , wr_623  , wr_618  );
  not  g591( wr_625  ,           wr_623  );
  nor  g592( wr_634  , wr_633  , wr_628  );
  not  g593( wr_635  ,           wr_633  );
  nor  g594( wr_644  , wr_643  , wr_638  );
  not  g595( wr_645  ,           wr_643  );
  nor  g596( wr_654  , wr_653  , wr_648  );
  not  g597( wr_655  ,           wr_653  );
  nor  g598( wr_669  , wr_543  , wr_668  );
  not  g599( wr_670  ,           wr_543  );
  nor  g600( wr_721  , wr_158  , wr_156  );
  nor  g601( wr_730  , wr_643  , G3705   );
  nor  g602( wr_252  , wr_249  , G2247   );
  nor  g603( wr_256  , wr_241  , G2253   );
  nor  g604( wr_281  , wr_259  , G2239   );
  nor  g605( wr_294  , wr_291  , G2236   );
  nor  g606( wr_447  , wr_446  , wr_441  );
  nor  g607( wr_452  , wr_436  , wr_451  );
  nor  g608( wr_480  , wr_460  , wr_479  );
  nor  g609( wr_496  , wr_495  , wr_490  );
  nor  g610( wr_578  , wr_577  , wr_572  );
  nor  g611( wr_588  , wr_587  , wr_582  );
  nor  g612( wr_608  , wr_607  , wr_602  );
  nor  g613( wr_694  , wr_577  , G3729   );
  not  g614( wr_236  ,           wr_235  );
  not  g615( wr_429  ,           wr_427  );
  nor  g616( wr_461  , wr_460  , G4420   );
  nor  g617( wr_238  , wr_235  , G2256   );
  nor  g618( wr_315  , wr_314  , G2224   );
  nor  g619( wr_349  , wr_330  , G2218   );
  nor  g620( wr_428  , wr_427  , wr_422  );
  nor  g621( wr_519  , wr_518  , G4405   );
  nor  g622( wr_553  , wr_534  , G4400   );
  nor  g623( wr_701  , wr_607  , G3737   );
  nor  g624( wr_716  , wr_633  , G3711   );
  nor  g625( wr_468  , wr_446  , G4427   );
  not  g626( wr_599  ,           wr_597  );
  not  g627( wr_1320 ,           wr_1319 );
  not  g628( wr_1322 ,           wr_1315 );
  nor  g629( wr_598  , wr_597  , wr_592  );
  nor  g630( wr_1389 , wr_1284 , wr_1283 );
  not  g631( wr_1308 ,           wr_1307 );
  not  g632( wr_1310 ,           wr_1303 );
  nor  g633( wr_437  , wr_436  , G4432   );
  nor  g634( wr_690  , wr_587  , G3743   );
  nor  g635( wr_1398 , wr_1276 , wr_1272 );
  nor  g636( wr_2545 , wr_259  , wr_279  );
  nor  g637( wr_2963 , wr_190  , wr_184  );
  nor  g638( wr_3283 , wr_159  , wr_155  );
  not  g639( wr_905  ,           wr_904  );
  not  g640( wr_910  ,           wr_909  );
  not  g641( wr_925  ,           wr_920  );
  not  g642( wr_927  ,           wr_916  );
  not  g643( wr_1131 ,           wr_1130 );
  not  g644( wr_1133 ,           wr_1126 );
  not  g645( wr_1147 ,           wr_1142 );
  not  g646( wr_1149 ,           wr_1138 );
  not  g647( wr_1259 ,           wr_1258 );
  not  g648( wr_1261 ,           wr_1254 );
  not  g649( wr_1277 ,           wr_1276 );
  not  g650( wr_1279 ,           wr_1272 );
  not  g651( wr_1296 ,           wr_1295 );
  not  g652( wr_1298 ,           wr_1291 );
  not  g653( wr_219  ,           wr_218  );
  nor  g654( wr_301  , wr_300  , G2230   );
  nor  g655( wr_505  , wr_504  , G4410   );
  nor  g656( wr_693  , wr_597  , G3749   );
  nor  g657( wr_712  , wr_623  , G3717   );
  nor  g658( wr_715  , wr_653  , G3723   );
  not  g659( wr_801  ,           wr_800  );
  not  g660( wr_806  ,           wr_805  );
  not  g661( wr_812  ,           wr_811  );
  not  g662( wr_817  ,           wr_816  );
  nor  g663( wr_912  , wr_909  , wr_904  );
  nor  g664( wr_966  , wr_965  , wr_961  );
  nor  g665( wr_1362 , wr_1234 , wr_1230 );
  nor  g666( wr_221  , wr_218  , G1486   );
  nor  g667( wr_808  , wr_805  , wr_800  );
  nor  g668( wr_819  , wr_816  , wr_811  );
  not  g669( wr_833  ,           wr_832  );
  not  g670( wr_838  ,           wr_837  );
  not  g671( wr_844  ,           wr_843  );
  not  g672( wr_864  ,           wr_848  );
  not  g673( wr_942  ,           wr_936  );
  not  g674( wr_944  ,           wr_932  );
  not  g675( wr_1055 ,           wr_1054 );
  not  g676( wr_1057 ,           wr_1050 );
  not  g677( wr_1083 ,           wr_1066 );
  not  g678( wr_1085 ,           wr_1062 );
  not  g679( wr_1164 ,           wr_1158 );
  not  g680( wr_1166 ,           wr_1154 );
  not  g681( wr_1178 ,           wr_1171 );
  nor  g682( wr_1188 , wr_1187 , wr_1183 );
  not  g683( wr_1223 ,           wr_1222 );
  not  g684( wr_1225 ,           wr_1218 );
  not  g685( wr_1338 ,           wr_1183 );
  not  g686( wr_1754 ,           wr_1753 );
  not  g687( wr_1761 ,           wr_1759 );
  not  g688( wr_1812 ,           wr_1810 );
  not  g689( wr_2169 ,           wr_2168 );
  not  g690( wr_2174 ,           wr_2172 );
  not  g691( wr_2223 ,           wr_2221 );
  not  g692( wr_790  ,           wr_789  );
  not  g693( wr_795  ,           wr_794  );
  nor  g694( wr_840  , wr_837  , wr_832  );
  nor  g695( wr_866  , wr_848  , wr_843  );
  nor  g696( wr_975  , wr_953  , wr_949  );
  nor  g697( wr_1369 , wr_1222 , wr_1218 );
  nor  g698( wr_1384 , wr_1295 , wr_1291 );
  not  g699( wr_770  ,           wr_769  );
  nor  g700( wr_797  , wr_794  , wr_789  );
  not  g701( wr_870  ,           wr_869  );
  not  g702( wr_893  ,           wr_874  );
  not  g703( wr_954  ,           wr_953  );
  not  g704( wr_956  ,           wr_949  );
  not  g705( wr_1033 ,           wr_965  );
  not  g706( wr_1035 ,           wr_961  );
  not  g707( wr_1113 ,           wr_1094 );
  not  g708( wr_1115 ,           wr_1090 );
  not  g709( wr_1176 ,           wr_1175 );
  nor  g710( wr_1197 , wr_1175 , wr_1171 );
  not  g711( wr_1247 ,           wr_1246 );
  not  g712( wr_1249 ,           wr_1242 );
  not  g713( wr_1336 ,           wr_1187 );
  not  g714( wr_1972 ,           wr_1971 );
  not  g715( wr_1974 ,           wr_1967 );
  not  g716( wr_2024 ,           wr_2022 );
  nor  g717( wr_440  , wr_427  , G4437   );
  nor  g718( wr_508  , wr_495  , G4415   );
  not  g719( wr_783  ,           wr_782  );
  nor  g720( wr_895  , wr_874  , wr_869  );
  not  g721( wr_775  ,           wr_774  );
  nor  g722( wr_786  , wr_782  , wr_785  );
  not  g723( wr_855  ,           wr_854  );
  not  g724( wr_860  ,           wr_859  );
  nor  g725( wr_1007 , wr_782  , wr_187  );
  not  g726( wr_1078 ,           wr_1077 );
  not  g727( wr_1080 ,           wr_1073 );
  nor  g728( wr_1095 , wr_1094 , wr_1090 );
  not  g729( wr_1235 ,           wr_1234 );
  not  g730( wr_1237 ,           wr_1230 );
  not  g731( wr_1663 ,           wr_1661 );
  nor  g732( wr_1707 , wr_1706 , wr_187  );
  not  g733( wr_1919 ,           wr_1917 );
  not  g734( wr_2078 ,           wr_2076 );
  nor  g735( wr_2123 , wr_2122 , wr_187  );
  nor  g736( wr_862  , wr_859  , wr_854  );
  nor  g737( wr_937  , wr_936  , wr_932  );
  nor  g738( wr_1653 , wr_300  , wr_291  );
  nor  g739( wr_2070 , wr_916  , wr_904  );
  nor  g740( wr_173  , wr_172  , wr_168  );
  nor  g741( wr_179  , wr_178  , wr_168  );
  nor  g742( wr_758  , wr_757  , wr_168  );
  nor  g743( wr_763  , wr_762  , wr_168  );
  nor  g744( wr_777  , wr_774  , wr_769  );
  nor  g745( wr_1102 , wr_1077 , wr_1073 );
  nor  g746( wr_1159 , wr_1158 , wr_1154 );
  not  g747( wr_1867 ,           wr_1865 );
  nor  g748( wr_1286 , wr_1285 , wr_1283 );
  nor  g749( wr_1358 , wr_1258 , wr_1254 );
  nor  g750( wr_1361 , wr_1246 , wr_1242 );
  nor  g751( wr_1380 , wr_1319 , wr_1315 );
  nor  g752( wr_1383 , wr_1307 , wr_1303 );
  not  g753( wr_1691 ,           wr_1690 );
  not  g754( wr_1695 ,           wr_1693 );
  not  g755( wr_2106 ,           wr_2105 );
  not  g756( wr_2110 ,           wr_2108 );
  nor  g757( wr_921  , wr_920  , wr_916  );
  not  g758( wr_1901 ,           wr_1900 );
  not  g759( wr_1903 ,           wr_1896 );
  nor  g760( wr_1067 , wr_1066 , wr_1062 );
  nor  g761( wr_1070 , wr_1054 , wr_1050 );
  nor  g762( wr_1143 , wr_1142 , wr_1138 );
  nor  g763( wr_1146 , wr_1130 , wr_1126 );
  nor  g764( wr_3009 , wr_172  , G38     );
  not  g765( wr_3002 ,           wr_3001 );
  nor  g766( wr_115  , wr_114  , wr_110  );
  nor  g767( wr_124  , wr_123  , wr_119  );
  not  g768( wr_368  ,           wr_367  );
  not  g769( wr_994  ,           wr_993  );
  nor  g770( wr_133  , wr_132  , wr_128  );
  nor  g771( wr_142  , wr_141  , wr_137  );
  nor  g772( wr_2571 , wr_172  , G38     );
  nor  g773( wr_151  , wr_150  , G5      );
  nor  g774( wr_162  , wr_161  , wr_160  );
  nor  g775( wr_192  , wr_191  , wr_184  );
  nor  g776( wr_199  , wr_198  , wr_195  );
  nor  g777( wr_206  , wr_205  , wr_202  );
  nor  g778( wr_213  , wr_212  , wr_209  );
  nor  g779( wr_308  , wr_307  , G2230   );
  nor  g780( wr_323  , wr_322  , G2224   );
  nor  g781( wr_333  , wr_332  , G2218   );
  not  g782( wr_341  ,           wr_340  );
  nor  g783( wr_381  , wr_191  , G1462   );
  nor  g784( wr_410  , wr_409  , G2211   );
  nor  g785( wr_512  , wr_511  , G4410   );
  nor  g786( wr_527  , wr_526  , G4405   );
  nor  g787( wr_537  , wr_536  , G4400   );
  not  g788( wr_545  ,           wr_544  );
  nor  g789( wr_626  , wr_625  , G3717   );
  nor  g790( wr_636  , wr_635  , G3711   );
  nor  g791( wr_646  , wr_645  , G3705   );
  nor  g792( wr_656  , wr_655  , G3723   );
  nor  g793( wr_671  , wr_670  , G4394   );
  not  g794( wr_722  ,           wr_721  );
  not  g795( wr_731  ,           wr_730  );
  nor  g796( wr_251  , wr_250  , wr_247  );
  nor  g797( wr_255  , wr_242  , wr_254  );
  nor  g798( wr_280  , wr_260  , wr_279  );
  nor  g799( wr_293  , wr_292  , wr_289  );
  nor  g800( wr_449  , wr_448  , G4427   );
  nor  g801( wr_454  , wr_453  , G4432   );
  nor  g802( wr_482  , wr_481  , G4420   );
  nor  g803( wr_498  , wr_497  , G4415   );
  nor  g804( wr_580  , wr_579  , G3729   );
  nor  g805( wr_590  , wr_589  , G3743   );
  nor  g806( wr_610  , wr_609  , G3737   );
  nor  g807( wr_261  , wr_260  , G2239   );
  not  g808( wr_695  ,           wr_694  );
  nor  g809( wr_237  , wr_236  , wr_233  );
  nor  g810( wr_376  , wr_205  , G106    );
  nor  g811( wr_390  , wr_212  , G1469   );
  nor  g812( wr_430  , wr_429  , G4437   );
  not  g813( wr_462  ,           wr_461  );
  nor  g814( wr_268  , wr_250  , G2247   );
  not  g815( wr_350  ,           wr_349  );
  not  g816( wr_554  ,           wr_553  );
  not  g817( wr_702  ,           wr_701  );
  not  g818( wr_717  ,           wr_716  );
  nor  g819( wr_600  , wr_599  , G3749   );
  nor  g820( wr_1321 , wr_1320 , wr_1315 );
  nor  g821( wr_1323 , wr_1319 , wr_1322 );
  not  g822( wr_1390 ,           wr_1389 );
  nor  g823( wr_243  , wr_242  , G2253   );
  nor  g824( wr_1309 , wr_1308 , wr_1303 );
  nor  g825( wr_1311 , wr_1307 , wr_1310 );
  nor  g826( wr_1626 , wr_579  , wr_572  );
  nor  g827( wr_2700 , wr_481  , wr_479  );
  nor  g828( wr_2785 , wr_409  , wr_407  );
  nor  g829( wr_3106 , wr_670  , wr_668  );
  not  g830( wr_316  ,           wr_315  );
  not  g831( wr_469  ,           wr_468  );
  not  g832( wr_520  ,           wr_519  );
  not  g833( wr_1399 ,           wr_1398 );
  not  g834( wr_2547 ,           wr_2545 );
  not  g835( wr_2966 ,           wr_2963 );
  not  g836( wr_3286 ,           wr_3283 );
  nor  g837( wr_372  , wr_198  , G1480   );
  nor  g838( wr_911  , wr_910  , wr_905  );
  nor  g839( wr_926  , wr_925  , wr_916  );
  nor  g840( wr_928  , wr_920  , wr_927  );
  nor  g841( wr_1132 , wr_1131 , wr_1126 );
  nor  g842( wr_1134 , wr_1130 , wr_1133 );
  nor  g843( wr_1148 , wr_1147 , wr_1138 );
  nor  g844( wr_1150 , wr_1142 , wr_1149 );
  nor  g845( wr_1260 , wr_1259 , wr_1254 );
  nor  g846( wr_1262 , wr_1258 , wr_1261 );
  nor  g847( wr_1278 , wr_1277 , wr_1272 );
  nor  g848( wr_1280 , wr_1276 , wr_1279 );
  nor  g849( wr_1297 , wr_1296 , wr_1291 );
  nor  g850( wr_1299 , wr_1295 , wr_1298 );
  nor  g851( wr_220  , wr_219  , wr_216  );
  not  g852( wr_691  ,           wr_690  );
  not  g853( wr_713  ,           wr_712  );
  nor  g854( wr_807  , wr_806  , wr_801  );
  nor  g855( wr_818  , wr_817  , wr_812  );
  not  g856( wr_967  ,           wr_966  );
  not  g857( wr_1363 ,           wr_1362 );
  nor  g858( wr_839  , wr_838  , wr_833  );
  nor  g859( wr_865  , wr_864  , wr_844  );
  nor  g860( wr_943  , wr_942  , wr_932  );
  nor  g861( wr_945  , wr_936  , wr_944  );
  nor  g862( wr_1056 , wr_1055 , wr_1050 );
  nor  g863( wr_1058 , wr_1054 , wr_1057 );
  nor  g864( wr_1084 , wr_1083 , wr_1062 );
  nor  g865( wr_1086 , wr_1066 , wr_1085 );
  nor  g866( wr_1165 , wr_1164 , wr_1154 );
  nor  g867( wr_1167 , wr_1158 , wr_1166 );
  not  g868( wr_1189 ,           wr_1188 );
  nor  g869( wr_1224 , wr_1223 , wr_1218 );
  nor  g870( wr_1226 , wr_1222 , wr_1225 );
  nor  g871( wr_1742 , wr_643  , wr_635  );
  nor  g872( wr_1743 , wr_645  , wr_633  );
  nor  g873( wr_1746 , wr_655  , wr_623  );
  nor  g874( wr_1747 , wr_653  , wr_625  );
  nor  g875( wr_1760 , wr_1759 , wr_1754 );
  nor  g876( wr_1762 , wr_1761 , wr_1753 );
  nor  g877( wr_1798 , wr_534  , wr_526  );
  nor  g878( wr_1799 , wr_536  , wr_518  );
  nor  g879( wr_1802 , wr_504  , wr_497  );
  nor  g880( wr_1803 , wr_511  , wr_495  );
  nor  g881( wr_1811 , wr_1810 , wr_670  );
  nor  g882( wr_1813 , wr_1812 , wr_543  );
  nor  g883( wr_2158 , wr_1298 , wr_1272 );
  nor  g884( wr_2159 , wr_1291 , wr_1279 );
  nor  g885( wr_2162 , wr_1315 , wr_1310 );
  nor  g886( wr_2163 , wr_1322 , wr_1303 );
  nor  g887( wr_2173 , wr_2172 , wr_2169 );
  nor  g888( wr_2175 , wr_2174 , wr_2168 );
  nor  g889( wr_2211 , wr_1171 , wr_1166 );
  nor  g890( wr_2212 , wr_1178 , wr_1154 );
  nor  g891( wr_2215 , wr_1138 , wr_1133 );
  nor  g892( wr_2216 , wr_1149 , wr_1126 );
  nor  g893( wr_2222 , wr_2221 , wr_1338 );
  nor  g894( wr_2224 , wr_2223 , wr_1183 );
  nor  g895( wr_796  , wr_795  , wr_790  );
  not  g896( wr_976  ,           wr_975  );
  not  g897( wr_1370 ,           wr_1369 );
  not  g898( wr_1385 ,           wr_1384 );
  nor  g899( wr_246  , wr_236  , G2256   );
  nor  g900( wr_304  , wr_292  , G2236   );
  nor  g901( wr_875  , wr_874  , wr_870  );
  nor  g902( wr_894  , wr_893  , wr_870  );
  nor  g903( wr_955  , wr_954  , wr_949  );
  nor  g904( wr_957  , wr_953  , wr_956  );
  nor  g905( wr_1034 , wr_1033 , wr_961  );
  nor  g906( wr_1036 , wr_965  , wr_1035 );
  nor  g907( wr_1114 , wr_1113 , wr_1090 );
  nor  g908( wr_1116 , wr_1094 , wr_1115 );
  not  g909( wr_1198 ,           wr_1197 );
  nor  g910( wr_1248 , wr_1247 , wr_1242 );
  nor  g911( wr_1250 , wr_1246 , wr_1249 );
  nor  g912( wr_1337 , wr_1336 , wr_1183 );
  nor  g913( wr_1339 , wr_1187 , wr_1338 );
  nor  g914( wr_1698 , wr_212  , wr_204  );
  nor  g915( wr_1699 , wr_211  , wr_205  );
  nor  g916( wr_1702 , wr_218  , wr_198  );
  nor  g917( wr_1703 , wr_219  , wr_197  );
  nor  g918( wr_1956 , wr_1296 , wr_1276 );
  nor  g919( wr_1957 , wr_1295 , wr_1277 );
  nor  g920( wr_1960 , wr_1319 , wr_1308 );
  nor  g921( wr_1961 , wr_1320 , wr_1307 );
  nor  g922( wr_1973 , wr_1972 , wr_1967 );
  nor  g923( wr_1975 , wr_1971 , wr_1974 );
  nor  g924( wr_2011 , wr_1175 , wr_1164 );
  nor  g925( wr_2012 , wr_1176 , wr_1158 );
  nor  g926( wr_2015 , wr_1142 , wr_1131 );
  nor  g927( wr_2016 , wr_1147 , wr_1130 );
  nor  g928( wr_2023 , wr_2022 , wr_1336 );
  nor  g929( wr_2025 , wr_2024 , wr_1187 );
  nor  g930( wr_2113 , wr_789  , wr_770  );
  nor  g931( wr_2114 , wr_790  , wr_769  );
  nor  g932( wr_2117 , wr_812  , wr_800  );
  nor  g933( wr_2118 , wr_811  , wr_801  );
  not  g934( wr_302  ,           wr_301  );
  not  g935( wr_438  ,           wr_437  );
  not  g936( wr_506  ,           wr_505  );
  nor  g937( wr_784  , wr_783  , wr_187  );
  nor  g938( wr_1177 , wr_1176 , wr_1171 );
  nor  g939( wr_1179 , wr_1175 , wr_1178 );
  nor  g940( wr_861  , wr_860  , wr_855  );
  nor  g941( wr_882  , wr_859  , wr_855  );
  not  g942( wr_1008 ,           wr_1007 );
  nor  g943( wr_1079 , wr_1078 , wr_1073 );
  nor  g944( wr_1081 , wr_1077 , wr_1080 );
  not  g945( wr_1096 ,           wr_1095 );
  nor  g946( wr_1236 , wr_1235 , wr_1230 );
  nor  g947( wr_1238 , wr_1234 , wr_1237 );
  nor  g948( wr_1649 , wr_330  , wr_322  );
  nor  g949( wr_1650 , wr_332  , wr_314  );
  nor  g950( wr_1654 , wr_307  , wr_292  );
  nor  g951( wr_1662 , wr_1661 , wr_409  );
  nor  g952( wr_1664 , wr_1663 , wr_339  );
  not  g953( wr_1711 ,           wr_1707 );
  nor  g954( wr_1731 , wr_609  , wr_577  );
  nor  g955( wr_1732 , wr_607  , wr_579  );
  nor  g956( wr_1734 , wr_599  , wr_587  );
  nor  g957( wr_1735 , wr_597  , wr_589  );
  nor  g958( wr_1787 , wr_460  , wr_448  );
  nor  g959( wr_1788 , wr_481  , wr_446  );
  nor  g960( wr_1790 , wr_436  , wr_429  );
  nor  g961( wr_1791 , wr_453  , wr_427  );
  nor  g962( wr_1906 , wr_795  , wr_774  );
  nor  g963( wr_1907 , wr_794  , wr_775  );
  nor  g964( wr_1910 , wr_816  , wr_806  );
  nor  g965( wr_1911 , wr_817  , wr_805  );
  nor  g966( wr_1918 , wr_1917 , wr_783  );
  nor  g967( wr_1920 , wr_1919 , wr_782  );
  nor  g968( wr_2066 , wr_949  , wr_944  );
  nor  g969( wr_2067 , wr_956  , wr_932  );
  nor  g970( wr_2071 , wr_927  , wr_905  );
  nor  g971( wr_2077 , wr_2076 , wr_1035 );
  nor  g972( wr_2079 , wr_2078 , wr_961  );
  not  g973( wr_2127 ,           wr_2123 );
  nor  g974( wr_2147 , wr_1230 , wr_1225 );
  nor  g975( wr_2148 , wr_1237 , wr_1218 );
  nor  g976( wr_2150 , wr_1254 , wr_1249 );
  nor  g977( wr_2151 , wr_1261 , wr_1242 );
  nor  g978( wr_2200 , wr_1090 , wr_1080 );
  nor  g979( wr_2201 , wr_1115 , wr_1073 );
  nor  g980( wr_2203 , wr_1062 , wr_1057 );
  nor  g981( wr_2204 , wr_1085 , wr_1050 );
  nor  g982( wr_776  , wr_775  , wr_770  );
  not  g983( wr_938  ,           wr_937  );
  nor  g984( wr_1016 , wr_774  , wr_770  );
  nor  g985( wr_175  , wr_174  , wr_173  );
  nor  g986( wr_181  , wr_180  , wr_179  );
  nor  g987( wr_760  , wr_759  , wr_758  );
  nor  g988( wr_765  , wr_764  , wr_763  );
  not  g989( wr_1103 ,           wr_1102 );
  not  g990( wr_1160 ,           wr_1159 );
  nor  g991( wr_1854 , wr_953  , wr_942  );
  nor  g992( wr_1855 , wr_954  , wr_936  );
  nor  g993( wr_1858 , wr_920  , wr_910  );
  nor  g994( wr_1859 , wr_925  , wr_909  );
  nor  g995( wr_1866 , wr_1865 , wr_1033 );
  nor  g996( wr_1868 , wr_1867 , wr_965  );
  nor  g997( wr_1945 , wr_1234 , wr_1223 );
  nor  g998( wr_1946 , wr_1235 , wr_1222 );
  nor  g999( wr_1948 , wr_1258 , wr_1247 );
  nor g1000( wr_1949 , wr_1259 , wr_1246 );
  nor g1001( wr_2000 , wr_1094 , wr_1078 );
  nor g1002( wr_2001 , wr_1113 , wr_1077 );
  nor g1003( wr_2003 , wr_1066 , wr_1055 );
  nor g1004( wr_2004 , wr_1083 , wr_1054 );
  nor g1005( wr_1288 , wr_1287 , wr_1286 );
  not g1006( wr_1359 ,           wr_1358 );
  not g1007( wr_1381 ,           wr_1380 );
  nor g1008( wr_1638 , wr_260  , wr_249  );
  nor g1009( wr_1639 , wr_259  , wr_250  );
  nor g1010( wr_1641 , wr_242  , wr_235  );
  nor g1011( wr_1642 , wr_241  , wr_236  );
  nor g1012( wr_2055 , wr_870  , wr_854  );
  nor g1013( wr_2056 , wr_869  , wr_855  );
  nor g1014( wr_2058 , wr_844  , wr_832  );
  nor g1015( wr_2059 , wr_843  , wr_833  );
  nor g1016( wr_1002 , wr_794  , wr_790  );
  nor g1017( wr_1694 , wr_1693 , wr_1691 );
  nor g1018( wr_1696 , wr_1695 , wr_1690 );
  nor g1019( wr_2109 , wr_2108 , wr_2106 );
  nor g1020( wr_2111 , wr_2110 , wr_2105 );
  nor g1021( wr_375  , wr_219  , G1486   );
  nor g1022( wr_849  , wr_848  , wr_844  );
  nor g1023( wr_852  , wr_837  , wr_833  );
  nor g1024( wr_924  , wr_909  , wr_905  );
  nor g1025( wr_1843 , wr_874  , wr_860  );
  nor g1026( wr_1844 , wr_893  , wr_859  );
  nor g1027( wr_1846 , wr_848  , wr_838  );
  nor g1028( wr_1847 , wr_864  , wr_837  );
  not g1029( wr_922  ,           wr_921  );
  nor g1030( wr_1902 , wr_1901 , wr_1896 );
  nor g1031( wr_1904 , wr_1900 , wr_1903 );
  not g1032( wr_1068 ,           wr_1067 );
  not g1033( wr_1144 ,           wr_1143 );
  not g1034( wr_3010 ,           wr_3009 );
  nor g1035( wr_998  , wr_816  , wr_812  );
  nor g1036( wr_1001 , wr_805  , wr_801  );
  not g1037( wr_116  ,           wr_115  );
  not g1038( wr_125  ,           wr_124  );
  not g1039( wr_134  ,           wr_133  );
  not g1040( wr_143  ,           wr_142  );
  not g1041( wr_2573 ,           wr_2571 );
  not g1042( G292    ,           wr_151  );
  not g1043( G281    ,           wr_151  );
  nor g1044( wr_194  , wr_193  , wr_192  );
  nor g1045( wr_215  , wr_214  , wr_213  );
  nor g1046( wr_334  , wr_333  , wr_331  );
  not g1047( wr_382  ,           wr_381  );
  nor g1048( wr_411  , wr_410  , wr_408  );
  nor g1049( wr_538  , wr_537  , wr_535  );
  nor g1050( wr_627  , wr_626  , wr_624  );
  nor g1051( wr_647  , wr_646  , wr_644  );
  nor g1052( wr_657  , wr_656  , wr_654  );
  nor g1053( wr_672  , wr_671  , wr_669  );
  nor g1054( wr_201  , wr_200  , wr_199  );
  nor g1055( wr_208  , wr_207  , wr_206  );
  nor g1056( wr_309  , wr_308  , wr_306  );
  nor g1057( wr_324  , wr_323  , wr_321  );
  nor g1058( wr_513  , wr_512  , wr_510  );
  nor g1059( wr_528  , wr_527  , wr_525  );
  nor g1060( wr_637  , wr_636  , wr_634  );
  nor g1061( wr_253  , wr_252  , wr_251  );
  nor g1062( wr_257  , wr_256  , wr_255  );
  nor g1063( wr_282  , wr_281  , wr_280  );
  nor g1064( wr_295  , wr_294  , wr_293  );
  nor g1065( wr_450  , wr_449  , wr_447  );
  nor g1066( wr_455  , wr_454  , wr_452  );
  nor g1067( wr_483  , wr_482  , wr_480  );
  nor g1068( wr_499  , wr_498  , wr_496  );
  nor g1069( wr_581  , wr_580  , wr_578  );
  nor g1070( wr_591  , wr_590  , wr_588  );
  nor g1071( wr_611  , wr_610  , wr_608  );
  not g1072( wr_262  ,           wr_261  );
  nor g1073( wr_239  , wr_238  , wr_237  );
  not g1074( wr_391  ,           wr_390  );
  nor g1075( wr_431  , wr_430  , wr_428  );
  nor g1076( wr_601  , wr_600  , wr_598  );
  nor g1077( wr_1324 , wr_1323 , wr_1321 );
  not g1078( wr_269  ,           wr_268  );
  nor g1079( wr_1312 , wr_1311 , wr_1309 );
  not g1080( wr_1628 ,           wr_1626 );
  not g1081( wr_2702 ,           wr_2700 );
  not g1082( wr_2788 ,           wr_2785 );
  not g1083( wr_3109 ,           wr_3106 );
  not g1084( wr_377  ,           wr_376  );
  nor g1085( wr_913  , wr_912  , wr_911  );
  nor g1086( wr_929  , wr_928  , wr_926  );
  nor g1087( wr_1135 , wr_1134 , wr_1132 );
  nor g1088( wr_1151 , wr_1150 , wr_1148 );
  nor g1089( wr_1263 , wr_1262 , wr_1260 );
  nor g1090( wr_1281 , wr_1280 , wr_1278 );
  nor g1091( wr_1300 , wr_1299 , wr_1297 );
  nor g1092( wr_222  , wr_221  , wr_220  );
  nor g1093( wr_809  , wr_808  , wr_807  );
  nor g1094( wr_820  , wr_819  , wr_818  );
  nor g1095( wr_841  , wr_840  , wr_839  );
  nor g1096( wr_867  , wr_866  , wr_865  );
  nor g1097( wr_946  , wr_945  , wr_943  );
  nor g1098( wr_1059 , wr_1058 , wr_1056 );
  nor g1099( wr_1087 , wr_1086 , wr_1084 );
  nor g1100( wr_1168 , wr_1167 , wr_1165 );
  nor g1101( wr_1227 , wr_1226 , wr_1224 );
  nor g1102( wr_1744 , wr_1743 , wr_1742 );
  nor g1103( wr_1748 , wr_1747 , wr_1746 );
  nor g1104( wr_1763 , wr_1762 , wr_1760 );
  nor g1105( wr_1800 , wr_1799 , wr_1798 );
  nor g1106( wr_1804 , wr_1803 , wr_1802 );
  nor g1107( wr_1814 , wr_1813 , wr_1811 );
  nor g1108( wr_2160 , wr_2159 , wr_2158 );
  nor g1109( wr_2164 , wr_2163 , wr_2162 );
  nor g1110( wr_2176 , wr_2175 , wr_2173 );
  nor g1111( wr_2213 , wr_2212 , wr_2211 );
  nor g1112( wr_2217 , wr_2216 , wr_2215 );
  nor g1113( wr_2225 , wr_2224 , wr_2222 );
  nor g1114( wr_798  , wr_797  , wr_796  );
  not g1115( wr_244  ,           wr_243  );
  not g1116( wr_876  ,           wr_875  );
  nor g1117( wr_896  , wr_895  , wr_894  );
  nor g1118( wr_958  , wr_957  , wr_955  );
  nor g1119( wr_1037 , wr_1036 , wr_1034 );
  nor g1120( wr_1117 , wr_1116 , wr_1114 );
  nor g1121( wr_1251 , wr_1250 , wr_1248 );
  nor g1122( wr_1340 , wr_1339 , wr_1337 );
  nor g1123( wr_1700 , wr_1699 , wr_1698 );
  nor g1124( wr_1704 , wr_1703 , wr_1702 );
  nor g1125( wr_1958 , wr_1957 , wr_1956 );
  nor g1126( wr_1962 , wr_1961 , wr_1960 );
  nor g1127( wr_1976 , wr_1975 , wr_1973 );
  nor g1128( wr_2013 , wr_2012 , wr_2011 );
  nor g1129( wr_2017 , wr_2016 , wr_2015 );
  nor g1130( wr_2026 , wr_2025 , wr_2023 );
  nor g1131( wr_2115 , wr_2114 , wr_2113 );
  nor g1132( wr_2119 , wr_2118 , wr_2117 );
  nor g1133( wr_787  , wr_786  , wr_784  );
  nor g1134( wr_1180 , wr_1179 , wr_1177 );
  not g1135( wr_165  ,           wr_162  );
  nor g1136( wr_863  , wr_862  , wr_861  );
  not g1137( wr_883  ,           wr_882  );
  nor g1138( wr_1082 , wr_1081 , wr_1079 );
  nor g1139( wr_1239 , wr_1238 , wr_1236 );
  nor g1140( wr_1651 , wr_1650 , wr_1649 );
  nor g1141( wr_1655 , wr_1654 , wr_1653 );
  nor g1142( wr_1665 , wr_1664 , wr_1662 );
  nor g1143( wr_1733 , wr_1732 , wr_1731 );
  nor g1144( wr_1736 , wr_1735 , wr_1734 );
  nor g1145( wr_1789 , wr_1788 , wr_1787 );
  nor g1146( wr_1792 , wr_1791 , wr_1790 );
  nor g1147( wr_1908 , wr_1907 , wr_1906 );
  nor g1148( wr_1912 , wr_1911 , wr_1910 );
  nor g1149( wr_1921 , wr_1920 , wr_1918 );
  nor g1150( wr_2068 , wr_2067 , wr_2066 );
  nor g1151( wr_2072 , wr_2071 , wr_2070 );
  nor g1152( wr_2080 , wr_2079 , wr_2077 );
  nor g1153( wr_2149 , wr_2148 , wr_2147 );
  nor g1154( wr_2152 , wr_2151 , wr_2150 );
  nor g1155( wr_2202 , wr_2201 , wr_2200 );
  nor g1156( wr_2205 , wr_2204 , wr_2203 );
  nor g1157( wr_778  , wr_777  , wr_776  );
  not g1158( wr_1017 ,           wr_1016 );
  nor g1159( wr_182  , wr_181  , wr_175  );
  nor g1160( wr_766  , wr_765  , wr_760  );
  nor g1161( wr_1856 , wr_1855 , wr_1854 );
  nor g1162( wr_1860 , wr_1859 , wr_1858 );
  nor g1163( wr_1869 , wr_1868 , wr_1866 );
  nor g1164( wr_1947 , wr_1946 , wr_1945 );
  nor g1165( wr_1950 , wr_1949 , wr_1948 );
  nor g1166( wr_2002 , wr_2001 , wr_2000 );
  nor g1167( wr_2005 , wr_2004 , wr_2003 );
  nor g1168( wr_1640 , wr_1639 , wr_1638 );
  nor g1169( wr_1643 , wr_1642 , wr_1641 );
  nor g1170( wr_2057 , wr_2056 , wr_2055 );
  nor g1171( wr_2060 , wr_2059 , wr_2058 );
  not g1172( wr_1003 ,           wr_1002 );
  nor g1173( wr_1697 , wr_1696 , wr_1694 );
  nor g1174( wr_2112 , wr_2111 , wr_2109 );
  not g1175( wr_373  ,           wr_372  );
  not g1176( wr_850  ,           wr_849  );
  nor g1177( wr_1845 , wr_1844 , wr_1843 );
  nor g1178( wr_1848 , wr_1847 , wr_1846 );
  nor g1179( wr_1905 , wr_1904 , wr_1902 );
  not g1180( wr_2567 ,           wr_181  );
  nor g1181( wr_3003 , wr_3002 , wr_181  );
  nor g1182( wr_3011 , wr_3010 , wr_181  );
  not g1183( wr_999  ,           wr_998  );
  nor g1184( wr_369  , wr_368  , wr_181  );
  nor g1185( wr_995  , wr_994  , wr_765  );
  nor g1186( wr_117  , wr_116  , wr_109  );
  nor g1187( wr_126  , wr_125  , wr_118  );
  nor g1188( wr_135  , wr_134  , wr_127  );
  nor g1189( wr_144  , wr_143  , wr_136  );
  nor g1190( wr_1564 , wr_162  , wr_164  );
  nor g1191( wr_2572 , wr_2571 , wr_181  );
  nor g1192( wr_2566 , wr_367  , wr_181  );
  not g1193( wr_2580 ,           wr_175  );
  nor g1194( wr_163  , wr_162  , G4526   );
  nor g1195( wr_723  , wr_722  , wr_627  );
  nor g1196( wr_1540 , wr_722  , wr_647  );
  nor g1197( wr_2380 , wr_341  , wr_334  );
  nor g1198( wr_2442 , wr_382  , wr_215  );
  nor g1199( wr_2614 , wr_545  , wr_538  );
  nor g1200( wr_2776 , wr_411  , wr_334  );
  nor g1201( wr_2954 , wr_215  , wr_194  );
  nor g1202( wr_3097 , wr_672  , wr_538  );
  nor g1203( wr_3274 , wr_647  , wr_162  );
  nor g1204( wr_732  , wr_731  , wr_627  );
  nor g1205( wr_342  , wr_341  , wr_309  );
  nor g1206( wr_383  , wr_382  , wr_201  );
  nor g1207( wr_546  , wr_545  , wr_513  );
  nor g1208( wr_1512 , wr_647  , wr_627  );
  nor g1209( wr_2352 , wr_334  , wr_309  );
  nor g1210( wr_2414 , wr_215  , wr_201  );
  nor g1211( wr_2586 , wr_538  , wr_513  );
  nor g1212( wr_412  , wr_334  , wr_295  );
  nor g1213( wr_673  , wr_538  , wr_499  );
  nor g1214( wr_696  , wr_695  , wr_591  );
  nor g1215( wr_1585 , wr_591  , wr_581  );
  nor g1216( wr_1588 , wr_611  , wr_591  );
  nor g1217( wr_2504 , wr_282  , wr_257  );
  nor g1218( wr_2507 , wr_257  , wr_253  );
  nor g1219( wr_2659 , wr_483  , wr_455  );
  nor g1220( wr_2662 , wr_455  , wr_450  );
  nor g1221( wr_1602 , wr_695  , wr_611  );
  nor g1222( wr_2521 , wr_262  , wr_253  );
  nor g1223( wr_2676 , wr_462  , wr_450  );
  nor g1224( wr_283  , wr_253  , wr_239  );
  nor g1225( wr_351  , wr_350  , wr_309  );
  nor g1226( wr_484  , wr_450  , wr_431  );
  nor g1227( wr_555  , wr_554  , wr_513  );
  nor g1228( wr_703  , wr_702  , wr_591  );
  nor g1229( wr_718  , wr_717  , wr_627  );
  nor g1230( wr_1509 , wr_637  , wr_627  );
  nor g1231( wr_1534 , wr_731  , wr_637  );
  nor g1232( wr_2349 , wr_324  , wr_309  );
  nor g1233( wr_2374 , wr_350  , wr_324  );
  nor g1234( wr_2411 , wr_208  , wr_201  );
  nor g1235( wr_2436 , wr_391  , wr_208  );
  nor g1236( wr_2583 , wr_528  , wr_513  );
  nor g1237( wr_2608 , wr_554  , wr_528  );
  nor g1238( wr_1443 , wr_309  , wr_295  );
  nor g1239( wr_1480 , wr_513  , wr_499  );
  nor g1240( wr_1611 , wr_611  , wr_581  );
  nor g1241( wr_2530 , wr_282  , wr_253  );
  nor g1242( wr_2685 , wr_483  , wr_450  );
  nor g1243( wr_263  , wr_262  , wr_257  );
  nor g1244( wr_463  , wr_462  , wr_455  );
  nor g1245( wr_612  , wr_611  , wr_601  );
  nor g1246( wr_658  , wr_657  , wr_647  );
  nor g1247( wr_1391 , wr_1390 , wr_1324 );
  nor g1248( wr_1434 , wr_257  , wr_239  );
  nor g1249( wr_1453 , wr_455  , wr_431  );
  nor g1250( wr_270  , wr_269  , wr_257  );
  nor g1251( wr_317  , wr_316  , wr_309  );
  nor g1252( wr_470  , wr_469  , wr_455  );
  nor g1253( wr_521  , wr_520  , wr_513  );
  nor g1254( wr_1400 , wr_1399 , wr_1324 );
  nor g1255( wr_1464 , wr_601  , wr_591  );
  nor g1256( wr_1470 , wr_657  , wr_627  );
  nor g1257( wr_378  , wr_377  , wr_201  );
  nor g1258( wr_692  , wr_691  , wr_601  );
  nor g1259( wr_714  , wr_713  , wr_657  );
  nor g1260( wr_968  , wr_967  , wr_929  );
  nor g1261( wr_1038 , wr_929  , wr_913  );
  nor g1262( wr_1341 , wr_1151 , wr_1135 );
  nor g1263( wr_1364 , wr_1363 , wr_1263 );
  nor g1264( wr_223  , wr_222  , wr_215  );
  nor g1265( wr_821  , wr_820  , wr_809  );
  nor g1266( wr_1190 , wr_1189 , wr_1151 );
  nor g1267( wr_1424 , wr_222  , wr_201  );
  nor g1268( wr_392  , wr_391  , wr_201  );
  nor g1269( wr_897  , wr_867  , wr_841  );
  nor g1270( wr_977  , wr_976  , wr_929  );
  nor g1271( wr_1118 , wr_1087 , wr_1059 );
  nor g1272( wr_1371 , wr_1370 , wr_1263 );
  nor g1273( wr_1386 , wr_1385 , wr_1324 );
  not g1274( wr_1745 ,           wr_1744 );
  not g1275( wr_1749 ,           wr_1748 );
  not g1276( wr_1767 ,           wr_1763 );
  not g1277( wr_1801 ,           wr_1800 );
  not g1278( wr_1805 ,           wr_1804 );
  not g1279( wr_1818 ,           wr_1814 );
  not g1280( wr_2161 ,           wr_2160 );
  not g1281( wr_2165 ,           wr_2164 );
  not g1282( wr_2180 ,           wr_2176 );
  not g1283( wr_2214 ,           wr_2213 );
  not g1284( wr_2218 ,           wr_2217 );
  not g1285( wr_2229 ,           wr_2225 );
  nor g1286( wr_1199 , wr_1198 , wr_1151 );
  not g1287( wr_1635 ,           wr_581  );
  nor g1288( wr_1776 , wr_1748 , wr_1744 );
  nor g1289( wr_1827 , wr_1804 , wr_1800 );
  nor g1290( wr_2189 , wr_2164 , wr_2160 );
  nor g1291( wr_2238 , wr_2217 , wr_2213 );
  not g1292( wr_2554 ,           wr_282  );
  not g1293( wr_2709 ,           wr_483  );
  nor g1294( wr_245  , wr_244  , wr_239  );
  nor g1295( wr_303  , wr_302  , wr_295  );
  nor g1296( wr_439  , wr_438  , wr_431  );
  nor g1297( wr_507  , wr_506  , wr_499  );
  nor g1298( wr_877  , wr_876  , wr_867  );
  nor g1299( wr_1264 , wr_1263 , wr_1251 );
  nor g1300( wr_1325 , wr_1324 , wr_1312 );
  not g1301( wr_1701 ,           wr_1700 );
  not g1302( wr_1705 ,           wr_1704 );
  not g1303( wr_1959 ,           wr_1958 );
  not g1304( wr_1963 ,           wr_1962 );
  not g1305( wr_1980 ,           wr_1976 );
  not g1306( wr_2014 ,           wr_2013 );
  not g1307( wr_2018 ,           wr_2017 );
  not g1308( wr_2030 ,           wr_2026 );
  not g1309( wr_2116 ,           wr_2115 );
  not g1310( wr_2120 ,           wr_2119 );
  nor g1311( wr_1009 , wr_1008 , wr_820  );
  nor g1312( wr_1097 , wr_1096 , wr_1087 );
  nor g1313( wr_1720 , wr_1704 , wr_1700 );
  nor g1314( wr_1989 , wr_1962 , wr_1958 );
  nor g1315( wr_2039 , wr_2017 , wr_2013 );
  nor g1316( wr_2136 , wr_2119 , wr_2115 );
  not g1317( wr_2287 ,           wr_411  );
  not g1318( wr_2307 ,           wr_194  );
  not g1319( wr_2563 ,           wr_672  );
  nor g1320( wr_884  , wr_883  , wr_867  );
  nor g1321( wr_939  , wr_938  , wr_929  );
  not g1322( wr_1622 ,           wr_611  );
  not g1323( wr_1652 ,           wr_1651 );
  not g1324( wr_1656 ,           wr_1655 );
  not g1325( wr_1669 ,           wr_1665 );
  not g1326( wr_1737 ,           wr_1736 );
  not g1327( wr_1739 ,           wr_1733 );
  not g1328( wr_1793 ,           wr_1792 );
  not g1329( wr_1795 ,           wr_1789 );
  not g1330( wr_1909 ,           wr_1908 );
  not g1331( wr_1913 ,           wr_1912 );
  not g1332( wr_1925 ,           wr_1921 );
  not g1333( wr_2069 ,           wr_2068 );
  not g1334( wr_2073 ,           wr_2072 );
  not g1335( wr_2084 ,           wr_2080 );
  not g1336( wr_2153 ,           wr_2152 );
  not g1337( wr_2155 ,           wr_2149 );
  not g1338( wr_2206 ,           wr_2205 );
  not g1339( wr_2208 ,           wr_2202 );
  not g1340( wr_2541 ,           wr_253  );
  not g1341( wr_2696 ,           wr_450  );
  nor g1342( wr_1018 , wr_1017 , wr_820  );
  nor g1343( wr_1104 , wr_1103 , wr_1087 );
  nor g1344( wr_1161 , wr_1160 , wr_1151 );
  nor g1345( wr_1678 , wr_1655 , wr_1651 );
  nor g1346( wr_1934 , wr_1912 , wr_1908 );
  nor g1347( wr_2093 , wr_2072 , wr_2068 );
  not g1348( wr_183  ,           wr_182  );
  not g1349( wr_767  ,           wr_766  );
  nor g1350( wr_1360 , wr_1359 , wr_1251 );
  nor g1351( wr_1382 , wr_1381 , wr_1312 );
  not g1352( wr_1568 ,           wr_647  );
  not g1353( wr_1857 ,           wr_1856 );
  not g1354( wr_1861 ,           wr_1860 );
  not g1355( wr_1873 ,           wr_1869 );
  not g1356( wr_1951 ,           wr_1950 );
  not g1357( wr_1953 ,           wr_1947 );
  not g1358( wr_2006 ,           wr_2005 );
  not g1359( wr_2008 ,           wr_2002 );
  not g1360( wr_2408 ,           wr_334  );
  not g1361( wr_2470 ,           wr_215  );
  not g1362( wr_2642 ,           wr_538  );
  not g1363( wr_1575 ,           wr_601  );
  nor g1364( wr_1882 , wr_1860 , wr_1856 );
  not g1365( wr_2494 ,           wr_239  );
  not g1366( wr_2649 ,           wr_431  );
  not g1367( wr_1644 ,           wr_1643 );
  not g1368( wr_1646 ,           wr_1640 );
  not g1369( wr_2061 ,           wr_2060 );
  not g1370( wr_2063 ,           wr_2057 );
  nor g1371( wr_1004 , wr_1003 , wr_820  );
  not g1372( wr_1531 ,           wr_657  );
  not g1373( wr_1728 ,           wr_1697 );
  not g1374( wr_2144 ,           wr_2112 );
  not g1375( wr_2371 ,           wr_295  );
  not g1376( wr_2433 ,           wr_222  );
  not g1377( wr_2605 ,           wr_499  );
  nor g1378( wr_374  , wr_373  , wr_222  );
  nor g1379( wr_851  , wr_850  , wr_841  );
  nor g1380( wr_923  , wr_922  , wr_913  );
  nor g1381( wr_1535 , wr_647  , wr_637  );
  not g1382( wr_1605 ,           wr_591  );
  not g1383( wr_1849 ,           wr_1848 );
  not g1384( wr_1851 ,           wr_1845 );
  nor g1385( wr_2375 , wr_334  , wr_324  );
  nor g1386( wr_2437 , wr_215  , wr_208  );
  not g1387( wr_2524 ,           wr_257  );
  nor g1388( wr_2609 , wr_538  , wr_528  );
  not g1389( wr_2679 ,           wr_455  );
  nor g1390( wr_1069 , wr_1068 , wr_1059 );
  nor g1391( wr_1145 , wr_1144 , wr_1135 );
  not g1392( wr_1942 ,           wr_1905 );
  nor g1393( wr_3004 , wr_3001 , wr_2567 );
  nor g1394( wr_3012 , wr_3009 , wr_2567 );
  not g1395( wr_1561 ,           wr_637  );
  not g1396( wr_2401 ,           wr_324  );
  not g1397( wr_2463 ,           wr_208  );
  not g1398( wr_2635 ,           wr_528  );
  nor g1399( wr_1553 , wr_647  , wr_164  );
  nor g1400( wr_1000 , wr_999  , wr_809  );
  not g1401( wr_1550 ,           wr_627  );
  not g1402( wr_2390 ,           wr_309  );
  not g1403( wr_2452 ,           wr_201  );
  not g1404( wr_2624 ,           wr_513  );
  nor g1405( wr_370  , wr_369  , wr_366  );
  nor g1406( wr_996  , wr_995  , wr_992  );
  not g1407( G404    ,           wr_117  );
  not g1408( G406    ,           wr_126  );
  nor g1409( wr_1627 , wr_1626 , wr_611  );
  nor g1410( wr_2546 , wr_2545 , wr_253  );
  nor g1411( wr_2574 , wr_2573 , wr_2567 );
  nor g1412( wr_2701 , wr_2700 , wr_450  );
  not g1413( G408    ,           wr_135  );
  not g1414( G410    ,           wr_144  );
  nor g1415( wr_1565 , wr_1564 , wr_721  );
  nor g1416( wr_1621 , wr_694  , wr_611  );
  nor g1417( wr_2540 , wr_261  , wr_253  );
  nor g1418( wr_2568 , wr_368  , wr_2567 );
  nor g1419( wr_2695 , wr_461  , wr_450  );
  nor g1420( wr_166  , wr_165  , wr_164  );
  not g1421( wr_724  ,           wr_723  );
  not g1422( wr_1541 ,           wr_1540 );
  not g1423( wr_2381 ,           wr_2380 );
  not g1424( wr_2443 ,           wr_2442 );
  not g1425( wr_2615 ,           wr_2614 );
  not g1426( wr_2778 ,           wr_2776 );
  not g1427( wr_2956 ,           wr_2954 );
  not g1428( wr_3099 ,           wr_3097 );
  not g1429( wr_3276 ,           wr_3274 );
  not g1430( wr_733  ,           wr_732  );
  not g1431( wr_343  ,           wr_342  );
  not g1432( wr_384  ,           wr_383  );
  not g1433( wr_547  ,           wr_546  );
  not g1434( wr_1513 ,           wr_1512 );
  not g1435( wr_2353 ,           wr_2352 );
  not g1436( wr_2415 ,           wr_2414 );
  not g1437( wr_2587 ,           wr_2586 );
  not g1438( wr_413  ,           wr_412  );
  not g1439( wr_674  ,           wr_673  );
  not g1440( wr_697  ,           wr_696  );
  not g1441( wr_1586 ,           wr_1585 );
  not g1442( wr_1589 ,           wr_1588 );
  not g1443( wr_2505 ,           wr_2504 );
  not g1444( wr_2508 ,           wr_2507 );
  not g1445( wr_2660 ,           wr_2659 );
  not g1446( wr_2663 ,           wr_2662 );
  nor g1447( wr_1603 , wr_1602 , wr_701  );
  nor g1448( wr_2522 , wr_2521 , wr_268  );
  nor g1449( wr_2677 , wr_2676 , wr_468  );
  not g1450( wr_284  ,           wr_283  );
  not g1451( wr_352  ,           wr_351  );
  not g1452( wr_485  ,           wr_484  );
  not g1453( wr_556  ,           wr_555  );
  not g1454( wr_704  ,           wr_703  );
  not g1455( wr_719  ,           wr_718  );
  not g1456( wr_1510 ,           wr_1509 );
  not g1457( wr_2350 ,           wr_2349 );
  not g1458( wr_2412 ,           wr_2411 );
  not g1459( wr_2584 ,           wr_2583 );
  not g1460( wr_1444 ,           wr_1443 );
  not g1461( wr_1481 ,           wr_1480 );
  not g1462( wr_264  ,           wr_263  );
  not g1463( wr_464  ,           wr_463  );
  not g1464( wr_613  ,           wr_612  );
  not g1465( wr_659  ,           wr_658  );
  not g1466( wr_1392 ,           wr_1391 );
  nor g1467( wr_2718 , wr_2380 , wr_349  );
  nor g1468( wr_2905 , wr_2442 , wr_390  );
  nor g1469( wr_3040 , wr_2614 , wr_553  );
  nor g1470( wr_3225 , wr_1540 , wr_730  );
  not g1471( wr_1435 ,           wr_1434 );
  not g1472( wr_1454 ,           wr_1453 );
  not g1473( wr_271  ,           wr_270  );
  not g1474( wr_318  ,           wr_317  );
  not g1475( wr_471  ,           wr_470  );
  not g1476( wr_522  ,           wr_521  );
  not g1477( wr_1401 ,           wr_1400 );
  not g1478( wr_1465 ,           wr_1464 );
  not g1479( wr_1471 ,           wr_1470 );
  not g1480( wr_969  ,           wr_968  );
  not g1481( wr_1039 ,           wr_1038 );
  not g1482( wr_1342 ,           wr_1341 );
  not g1483( wr_1365 ,           wr_1364 );
  not g1484( wr_224  ,           wr_223  );
  not g1485( wr_822  ,           wr_821  );
  not g1486( wr_1191 ,           wr_1190 );
  not g1487( wr_1425 ,           wr_1424 );
  not g1488( wr_393  ,           wr_392  );
  not g1489( wr_898  ,           wr_897  );
  not g1490( wr_978  ,           wr_977  );
  not g1491( wr_1119 ,           wr_1118 );
  not g1492( wr_1372 ,           wr_1371 );
  not g1493( wr_1387 ,           wr_1386 );
  nor g1494( wr_1764 , wr_1763 , wr_1749 );
  nor g1495( wr_1768 , wr_1748 , wr_1745 );
  nor g1496( wr_1773 , wr_1767 , wr_1749 );
  nor g1497( wr_1815 , wr_1814 , wr_1805 );
  nor g1498( wr_1819 , wr_1804 , wr_1801 );
  nor g1499( wr_1824 , wr_1818 , wr_1805 );
  nor g1500( wr_2177 , wr_2176 , wr_2165 );
  nor g1501( wr_2181 , wr_2164 , wr_2161 );
  nor g1502( wr_2186 , wr_2180 , wr_2165 );
  nor g1503( wr_2226 , wr_2225 , wr_2218 );
  nor g1504( wr_2230 , wr_2217 , wr_2214 );
  nor g1505( wr_2235 , wr_2229 , wr_2218 );
  not g1506( wr_1200 ,           wr_1199 );
  not g1507( wr_1777 ,           wr_1776 );
  not g1508( wr_1828 ,           wr_1827 );
  not g1509( wr_2190 ,           wr_2189 );
  not g1510( wr_2239 ,           wr_2238 );
  not g1511( wr_878  ,           wr_877  );
  not g1512( wr_1265 ,           wr_1264 );
  not g1513( wr_1326 ,           wr_1325 );
  nor g1514( wr_1708 , wr_1707 , wr_1705 );
  nor g1515( wr_1712 , wr_1704 , wr_1701 );
  nor g1516( wr_1717 , wr_1711 , wr_1705 );
  nor g1517( wr_1977 , wr_1976 , wr_1963 );
  nor g1518( wr_1981 , wr_1962 , wr_1959 );
  nor g1519( wr_1986 , wr_1980 , wr_1963 );
  nor g1520( wr_2027 , wr_2026 , wr_2018 );
  nor g1521( wr_2031 , wr_2017 , wr_2014 );
  nor g1522( wr_2036 , wr_2030 , wr_2018 );
  nor g1523( wr_2124 , wr_2123 , wr_2120 );
  nor g1524( wr_2128 , wr_2119 , wr_2116 );
  nor g1525( wr_2133 , wr_2127 , wr_2120 );
  not g1526( wr_1010 ,           wr_1009 );
  not g1527( wr_1098 ,           wr_1097 );
  not g1528( wr_1721 ,           wr_1720 );
  not g1529( wr_1990 ,           wr_1989 );
  not g1530( wr_2040 ,           wr_2039 );
  not g1531( wr_2137 ,           wr_2136 );
  not g1532( wr_379  ,           wr_378  );
  not g1533( wr_885  ,           wr_884  );
  not g1534( wr_940  ,           wr_939  );
  nor g1535( wr_1666 , wr_1665 , wr_1656 );
  nor g1536( wr_1670 , wr_1655 , wr_1652 );
  nor g1537( wr_1675 , wr_1669 , wr_1656 );
  nor g1538( wr_1738 , wr_1737 , wr_1733 );
  nor g1539( wr_1740 , wr_1736 , wr_1739 );
  nor g1540( wr_1794 , wr_1793 , wr_1789 );
  nor g1541( wr_1796 , wr_1792 , wr_1795 );
  nor g1542( wr_1922 , wr_1921 , wr_1913 );
  nor g1543( wr_1926 , wr_1912 , wr_1909 );
  nor g1544( wr_1931 , wr_1925 , wr_1913 );
  nor g1545( wr_2081 , wr_2080 , wr_2073 );
  nor g1546( wr_2085 , wr_2072 , wr_2069 );
  nor g1547( wr_2090 , wr_2084 , wr_2073 );
  nor g1548( wr_2154 , wr_2153 , wr_2149 );
  nor g1549( wr_2156 , wr_2152 , wr_2155 );
  nor g1550( wr_2207 , wr_2206 , wr_2202 );
  nor g1551( wr_2209 , wr_2205 , wr_2208 );
  not g1552( wr_1019 ,           wr_1018 );
  not g1553( wr_1105 ,           wr_1104 );
  not g1554( wr_1162 ,           wr_1161 );
  not g1555( wr_1679 ,           wr_1678 );
  not g1556( wr_1935 ,           wr_1934 );
  not g1557( wr_2094 ,           wr_2093 );
  nor g1558( wr_1870 , wr_1869 , wr_1861 );
  nor g1559( wr_1874 , wr_1860 , wr_1857 );
  nor g1560( wr_1879 , wr_1873 , wr_1861 );
  nor g1561( wr_1952 , wr_1951 , wr_1947 );
  nor g1562( wr_1954 , wr_1950 , wr_1953 );
  nor g1563( wr_2007 , wr_2006 , wr_2002 );
  nor g1564( wr_2009 , wr_2005 , wr_2008 );
  not g1565( wr_1883 ,           wr_1882 );
  nor g1566( wr_1645 , wr_1644 , wr_1640 );
  nor g1567( wr_1647 , wr_1643 , wr_1646 );
  nor g1568( wr_2062 , wr_2061 , wr_2057 );
  nor g1569( wr_2064 , wr_2060 , wr_2063 );
  not g1570( wr_1005 ,           wr_1004 );
  not g1571( wr_1536 ,           wr_1535 );
  nor g1572( wr_1850 , wr_1849 , wr_1845 );
  nor g1573( wr_1852 , wr_1848 , wr_1851 );
  not g1574( wr_2376 ,           wr_2375 );
  not g1575( wr_2438 ,           wr_2437 );
  not g1576( wr_2610 ,           wr_2609 );
  nor g1577( wr_3005 , wr_3004 , wr_3003 );
  nor g1578( wr_3013 , wr_3012 , wr_3011 );
  not g1579( wr_1554 ,           wr_1553 );
  nor g1580( wr_1612 , wr_1611 , wr_701  );
  nor g1581( wr_2531 , wr_2530 , wr_268  );
  nor g1582( wr_2686 , wr_2685 , wr_468  );
  not g1583( wr_371  ,           wr_370  );
  not g1584( wr_997  ,           wr_996  );
  nor g1585( wr_1629 , wr_1628 , wr_1622 );
  nor g1586( wr_2479 , G406    , G404    );
  nor g1587( wr_2548 , wr_2547 , wr_2541 );
  nor g1588( wr_2703 , wr_2702 , wr_2696 );
  nor g1589( wr_1623 , wr_695  , wr_1622 );
  nor g1590( wr_2542 , wr_262  , wr_2541 );
  nor g1591( wr_2575 , wr_2574 , wr_2572 );
  nor g1592( wr_2697 , wr_462  , wr_2696 );
  not g1593( wr_1566 ,           wr_1565 );
  nor g1594( wr_2473 , G410    , G408    );
  nor g1595( wr_2569 , wr_2568 , wr_2566 );
  nor g1596( wr_1569 , wr_1565 , wr_1568 );
  nor g1597( wr_167  , wr_166  , wr_163  );
  nor g1598( wr_725  , wr_724  , wr_657  );
  nor g1599( wr_1542 , wr_1541 , wr_637  );
  nor g1600( wr_2382 , wr_2381 , wr_324  );
  nor g1601( wr_2444 , wr_2443 , wr_208  );
  nor g1602( wr_2616 , wr_2615 , wr_528  );
  nor g1603( wr_2779 , wr_2778 , wr_324  );
  nor g1604( wr_2957 , wr_2956 , wr_208  );
  nor g1605( wr_3100 , wr_3099 , wr_528  );
  nor g1606( wr_3277 , wr_3276 , wr_637  );
  nor g1607( wr_734  , wr_733  , wr_637  );
  nor g1608( wr_1519 , wr_724  , wr_647  );
  nor g1609( wr_2359 , wr_343  , wr_334  );
  nor g1610( wr_2421 , wr_384  , wr_215  );
  nor g1611( wr_2593 , wr_547  , wr_538  );
  nor g1612( wr_2766 , wr_2353 , wr_411  );
  nor g1613( wr_2944 , wr_2415 , wr_194  );
  nor g1614( wr_3087 , wr_2587 , wr_672  );
  nor g1615( wr_3264 , wr_1513 , wr_162  );
  nor g1616( wr_344  , wr_343  , wr_295  );
  nor g1617( wr_414  , wr_413  , wr_324  );
  nor g1618( wr_548  , wr_547  , wr_499  );
  nor g1619( wr_675  , wr_674  , wr_528  );
  nor g1620( wr_698  , wr_697  , wr_611  );
  nor g1621( wr_1587 , wr_1586 , wr_611  );
  nor g1622( wr_1590 , wr_1589 , wr_695  );
  nor g1623( wr_2506 , wr_2505 , wr_253  );
  nor g1624( wr_2509 , wr_2508 , wr_262  );
  nor g1625( wr_2661 , wr_2660 , wr_450  );
  nor g1626( wr_2664 , wr_2663 , wr_462  );
  not g1627( wr_1606 ,           wr_1603 );
  not g1628( wr_2525 ,           wr_2522 );
  not g1629( wr_2680 ,           wr_2677 );
  nor g1630( wr_285  , wr_284  , wr_257  );
  nor g1631( wr_353  , wr_352  , wr_324  );
  nor g1632( wr_486  , wr_485  , wr_455  );
  nor g1633( wr_557  , wr_556  , wr_528  );
  nor g1634( wr_705  , wr_704  , wr_601  );
  nor g1635( wr_720  , wr_719  , wr_657  );
  nor g1636( wr_1511 , wr_1510 , wr_731  );
  nor g1637( wr_2351 , wr_2350 , wr_350  );
  nor g1638( wr_2413 , wr_2412 , wr_391  );
  nor g1639( wr_2585 , wr_2584 , wr_554  );
  nor g1640( wr_1445 , wr_1444 , wr_324  );
  nor g1641( wr_1482 , wr_1481 , wr_528  );
  nor g1642( wr_265  , wr_264  , wr_253  );
  nor g1643( wr_465  , wr_464  , wr_450  );
  nor g1644( wr_614  , wr_613  , wr_591  );
  nor g1645( wr_660  , wr_659  , wr_637  );
  nor g1646( wr_1393 , wr_1392 , wr_1312 );
  not g1647( wr_2719 ,           wr_2718 );
  nor g1648( wr_2856 , wr_2522 , wr_262  );
  not g1649( wr_2906 ,           wr_2905 );
  not g1650( wr_3041 ,           wr_3040 );
  nor g1651( wr_3177 , wr_2677 , wr_462  );
  not g1652( wr_3226 ,           wr_3225 );
  nor g1653( wr_3354 , wr_1603 , wr_695  );
  nor g1654( wr_1436 , wr_1435 , wr_282  );
  nor g1655( wr_1455 , wr_1454 , wr_483  );
  nor g1656( wr_272  , wr_271  , wr_239  );
  nor g1657( wr_319  , wr_318  , wr_295  );
  nor g1658( wr_472  , wr_471  , wr_431  );
  nor g1659( wr_523  , wr_522  , wr_499  );
  nor g1660( wr_1402 , wr_1401 , wr_1300 );
  nor g1661( wr_1466 , wr_1465 , wr_581  );
  nor g1662( wr_1472 , wr_1471 , wr_637  );
  nor g1663( wr_385  , wr_384  , wr_222  );
  nor g1664( wr_970  , wr_969  , wr_913  );
  nor g1665( wr_1040 , wr_1039 , wr_946  );
  nor g1666( wr_1343 , wr_1342 , wr_1168 );
  nor g1667( wr_1366 , wr_1365 , wr_1227 );
  nor g1668( wr_225  , wr_224  , wr_208  );
  nor g1669( wr_823  , wr_822  , wr_798  );
  nor g1670( wr_1192 , wr_1191 , wr_1135 );
  nor g1671( wr_1426 , wr_1425 , wr_208  );
  nor g1672( wr_394  , wr_393  , wr_208  );
  nor g1673( wr_899  , wr_898  , wr_896  );
  nor g1674( wr_979  , wr_978  , wr_946  );
  nor g1675( wr_1120 , wr_1119 , wr_1117 );
  nor g1676( wr_1373 , wr_1372 , wr_1251 );
  nor g1677( wr_1388 , wr_1387 , wr_1312 );
  not g1678( wr_1765 ,           wr_1764 );
  not g1679( wr_1769 ,           wr_1768 );
  not g1680( wr_1774 ,           wr_1773 );
  not g1681( wr_1816 ,           wr_1815 );
  not g1682( wr_1820 ,           wr_1819 );
  not g1683( wr_1825 ,           wr_1824 );
  not g1684( wr_2178 ,           wr_2177 );
  not g1685( wr_2182 ,           wr_2181 );
  not g1686( wr_2187 ,           wr_2186 );
  not g1687( wr_2227 ,           wr_2226 );
  not g1688( wr_2231 ,           wr_2230 );
  not g1689( wr_2236 ,           wr_2235 );
  nor g1690( wr_1201 , wr_1200 , wr_1168 );
  nor g1691( wr_1778 , wr_1777 , wr_1763 );
  nor g1692( wr_1829 , wr_1828 , wr_1814 );
  nor g1693( wr_2191 , wr_2190 , wr_2176 );
  nor g1694( wr_2240 , wr_2239 , wr_2225 );
  nor g1695( wr_879  , wr_878  , wr_863  );
  nor g1696( wr_1266 , wr_1265 , wr_1239 );
  nor g1697( wr_1327 , wr_1326 , wr_1300 );
  not g1698( wr_1709 ,           wr_1708 );
  not g1699( wr_1713 ,           wr_1712 );
  not g1700( wr_1718 ,           wr_1717 );
  not g1701( wr_1978 ,           wr_1977 );
  not g1702( wr_1982 ,           wr_1981 );
  not g1703( wr_1987 ,           wr_1986 );
  not g1704( wr_2028 ,           wr_2027 );
  not g1705( wr_2032 ,           wr_2031 );
  not g1706( wr_2037 ,           wr_2036 );
  not g1707( wr_2125 ,           wr_2124 );
  not g1708( wr_2129 ,           wr_2128 );
  not g1709( wr_2134 ,           wr_2133 );
  nor g1710( wr_1011 , wr_1010 , wr_809  );
  nor g1711( wr_1099 , wr_1098 , wr_1082 );
  nor g1712( wr_1722 , wr_1721 , wr_1707 );
  nor g1713( wr_1991 , wr_1990 , wr_1976 );
  nor g1714( wr_2041 , wr_2040 , wr_2026 );
  nor g1715( wr_2138 , wr_2137 , wr_2123 );
  nor g1716( wr_380  , wr_379  , wr_222  );
  nor g1717( wr_886  , wr_885  , wr_841  );
  nor g1718( wr_941  , wr_940  , wr_913  );
  not g1719( wr_1667 ,           wr_1666 );
  not g1720( wr_1671 ,           wr_1670 );
  not g1721( wr_1676 ,           wr_1675 );
  nor g1722( wr_1741 , wr_1740 , wr_1738 );
  nor g1723( wr_1797 , wr_1796 , wr_1794 );
  not g1724( wr_1923 ,           wr_1922 );
  not g1725( wr_1927 ,           wr_1926 );
  not g1726( wr_1932 ,           wr_1931 );
  not g1727( wr_2082 ,           wr_2081 );
  not g1728( wr_2086 ,           wr_2085 );
  not g1729( wr_2091 ,           wr_2090 );
  nor g1730( wr_2157 , wr_2156 , wr_2154 );
  nor g1731( wr_2210 , wr_2209 , wr_2207 );
  nor g1732( wr_1020 , wr_1019 , wr_798  );
  nor g1733( wr_1106 , wr_1105 , wr_1059 );
  nor g1734( wr_1163 , wr_1162 , wr_1135 );
  nor g1735( wr_1680 , wr_1679 , wr_1665 );
  nor g1736( wr_1936 , wr_1935 , wr_1921 );
  nor g1737( wr_2095 , wr_2094 , wr_2080 );
  nor g1738( wr_1514 , wr_1513 , wr_637  );
  not g1739( wr_1871 ,           wr_1870 );
  not g1740( wr_1875 ,           wr_1874 );
  not g1741( wr_1880 ,           wr_1879 );
  nor g1742( wr_1955 , wr_1954 , wr_1952 );
  nor g1743( wr_2010 , wr_2009 , wr_2007 );
  nor g1744( wr_2354 , wr_2353 , wr_324  );
  nor g1745( wr_2416 , wr_2415 , wr_208  );
  nor g1746( wr_2588 , wr_2587 , wr_528  );
  nor g1747( wr_1884 , wr_1883 , wr_1869 );
  nor g1748( wr_1648 , wr_1647 , wr_1645 );
  nor g1749( wr_2065 , wr_2064 , wr_2062 );
  nor g1750( wr_1006 , wr_1005 , wr_809  );
  nor g1751( wr_1537 , wr_1536 , wr_164  );
  nor g1752( wr_1853 , wr_1852 , wr_1850 );
  nor g1753( wr_1555 , wr_1554 , wr_162  );
  not g1754( wr_1613 ,           wr_1612 );
  not g1755( wr_2532 ,           wr_2531 );
  not g1756( wr_2687 ,           wr_2686 );
  nor g1757( wr_1604 , wr_1603 , wr_591  );
  nor g1758( wr_2523 , wr_2522 , wr_257  );
  nor g1759( wr_2678 , wr_2677 , wr_455  );
  nor g1760( wr_1630 , wr_1629 , wr_1627 );
  not g1761( wr_2480 ,           wr_2479 );
  nor g1762( wr_2549 , wr_2548 , wr_2546 );
  nor g1763( wr_2704 , wr_2703 , wr_2701 );
  nor g1764( wr_1624 , wr_1623 , wr_1621 );
  nor g1765( wr_2254 , wr_997  , wr_766  );
  nor g1766( wr_2326 , wr_371  , wr_182  );
  nor g1767( wr_2543 , wr_2542 , wr_2540 );
  not g1768( wr_2576 ,           wr_2575 );
  nor g1769( wr_2698 , wr_2697 , wr_2695 );
  nor g1770( wr_1567 , wr_1566 , wr_647  );
  not g1771( wr_2474 ,           wr_2473 );
  not g1772( G373    ,           wr_167  );
  not g1773( wr_726  ,           wr_725  );
  nor g1774( wr_2780 , wr_2779 , wr_2382 );
  nor g1775( wr_2958 , wr_2957 , wr_2444 );
  nor g1776( wr_3101 , wr_3100 , wr_2616 );
  nor g1777( wr_3278 , wr_3277 , wr_1542 );
  not g1778( wr_735  ,           wr_734  );
  nor g1779( wr_2720 , wr_2382 , wr_315  );
  nor g1780( wr_2907 , wr_2444 , wr_376  );
  nor g1781( wr_3042 , wr_2616 , wr_519  );
  nor g1782( wr_3227 , wr_1542 , wr_716  );
  not g1783( wr_1520 ,           wr_1519 );
  not g1784( wr_2360 ,           wr_2359 );
  not g1785( wr_2422 ,           wr_2421 );
  not g1786( wr_2594 ,           wr_2593 );
  not g1787( wr_2767 ,           wr_2766 );
  not g1788( wr_2945 ,           wr_2944 );
  not g1789( wr_3088 ,           wr_3087 );
  not g1790( wr_3265 ,           wr_3264 );
  not g1791( wr_345  ,           wr_344  );
  not g1792( wr_415  ,           wr_414  );
  not g1793( wr_549  ,           wr_548  );
  not g1794( wr_676  ,           wr_675  );
  not g1795( wr_699  ,           wr_698  );
  nor g1796( wr_1591 , wr_1590 , wr_1587 );
  nor g1797( wr_2510 , wr_2509 , wr_2506 );
  nor g1798( wr_2665 , wr_2664 , wr_2661 );
  nor g1799( wr_2823 , wr_2530 , wr_2525 );
  nor g1800( wr_3144 , wr_2685 , wr_2680 );
  nor g1801( wr_3321 , wr_1611 , wr_1606 );
  not g1802( wr_286  ,           wr_285  );
  not g1803( wr_354  ,           wr_353  );
  not g1804( wr_487  ,           wr_486  );
  not g1805( wr_558  ,           wr_557  );
  nor g1806( wr_2851 , wr_2509 , wr_243  );
  nor g1807( wr_3172 , wr_2664 , wr_437  );
  nor g1808( wr_3349 , wr_1590 , wr_690  );
  not g1809( wr_1446 ,           wr_1445 );
  not g1810( wr_1483 ,           wr_1482 );
  nor g1811( wr_2855 , wr_2525 , wr_261  );
  nor g1812( wr_3176 , wr_2680 , wr_461  );
  nor g1813( wr_3353 , wr_1606 , wr_694  );
  not g1814( wr_266  ,           wr_265  );
  not g1815( wr_466  ,           wr_465  );
  not g1816( wr_615  ,           wr_614  );
  not g1817( wr_661  ,           wr_660  );
  not g1818( wr_1394 ,           wr_1393 );
  nor g1819( wr_2777 , wr_2776 , wr_2719 );
  nor g1820( wr_2955 , wr_2954 , wr_2906 );
  nor g1821( wr_3098 , wr_3097 , wr_3041 );
  nor g1822( wr_3275 , wr_3274 , wr_3226 );
  not g1823( wr_1437 ,           wr_1436 );
  not g1824( wr_1456 ,           wr_1455 );
  not g1825( wr_1403 ,           wr_1402 );
  not g1826( wr_1467 ,           wr_1466 );
  not g1827( wr_1473 ,           wr_1472 );
  not g1828( wr_386  ,           wr_385  );
  not g1829( wr_971  ,           wr_970  );
  not g1830( wr_1041 ,           wr_1040 );
  not g1831( wr_1344 ,           wr_1343 );
  not g1832( wr_1367 ,           wr_1366 );
  not g1833( wr_226  ,           wr_225  );
  not g1834( wr_824  ,           wr_823  );
  not g1835( wr_1193 ,           wr_1192 );
  not g1836( wr_1427 ,           wr_1426 );
  not g1837( wr_395  ,           wr_394  );
  not g1838( wr_900  ,           wr_899  );
  not g1839( wr_980  ,           wr_979  );
  not g1840( wr_1121 ,           wr_1120 );
  nor g1841( wr_1766 , wr_1765 , wr_1745 );
  nor g1842( wr_1770 , wr_1769 , wr_1767 );
  nor g1843( wr_1775 , wr_1774 , wr_1744 );
  nor g1844( wr_1817 , wr_1816 , wr_1801 );
  nor g1845( wr_1821 , wr_1820 , wr_1818 );
  nor g1846( wr_1826 , wr_1825 , wr_1800 );
  nor g1847( wr_2179 , wr_2178 , wr_2161 );
  nor g1848( wr_2183 , wr_2182 , wr_2180 );
  nor g1849( wr_2188 , wr_2187 , wr_2160 );
  nor g1850( wr_2228 , wr_2227 , wr_2214 );
  nor g1851( wr_2232 , wr_2231 , wr_2229 );
  nor g1852( wr_2237 , wr_2236 , wr_2213 );
  not g1853( wr_1202 ,           wr_1201 );
  not g1854( wr_880  ,           wr_879  );
  not g1855( wr_1267 ,           wr_1266 );
  not g1856( wr_1328 ,           wr_1327 );
  nor g1857( wr_1710 , wr_1709 , wr_1701 );
  nor g1858( wr_1714 , wr_1713 , wr_1711 );
  nor g1859( wr_1719 , wr_1718 , wr_1700 );
  nor g1860( wr_1979 , wr_1978 , wr_1959 );
  nor g1861( wr_1983 , wr_1982 , wr_1980 );
  nor g1862( wr_1988 , wr_1987 , wr_1958 );
  nor g1863( wr_2029 , wr_2028 , wr_2014 );
  nor g1864( wr_2033 , wr_2032 , wr_2030 );
  nor g1865( wr_2038 , wr_2037 , wr_2013 );
  nor g1866( wr_2126 , wr_2125 , wr_2116 );
  nor g1867( wr_2130 , wr_2129 , wr_2127 );
  nor g1868( wr_2135 , wr_2134 , wr_2115 );
  not g1869( wr_1012 ,           wr_1011 );
  not g1870( wr_1100 ,           wr_1099 );
  nor g1871( wr_1668 , wr_1667 , wr_1652 );
  nor g1872( wr_1672 , wr_1671 , wr_1669 );
  nor g1873( wr_1677 , wr_1676 , wr_1651 );
  not g1874( wr_1784 ,           wr_1741 );
  not g1875( wr_1835 ,           wr_1797 );
  nor g1876( wr_1924 , wr_1923 , wr_1909 );
  nor g1877( wr_1928 , wr_1927 , wr_1925 );
  nor g1878( wr_1933 , wr_1932 , wr_1908 );
  nor g1879( wr_2083 , wr_2082 , wr_2069 );
  nor g1880( wr_2087 , wr_2086 , wr_2084 );
  nor g1881( wr_2092 , wr_2091 , wr_2068 );
  not g1882( wr_2197 ,           wr_2157 );
  not g1883( wr_2246 ,           wr_2210 );
  not g1884( wr_1021 ,           wr_1020 );
  not g1885( wr_1515 ,           wr_1514 );
  nor g1886( wr_1872 , wr_1871 , wr_1857 );
  nor g1887( wr_1876 , wr_1875 , wr_1873 );
  nor g1888( wr_1881 , wr_1880 , wr_1856 );
  not g1889( wr_1997 ,           wr_1955 );
  not g1890( wr_2047 ,           wr_2010 );
  not g1891( wr_2355 ,           wr_2354 );
  not g1892( wr_2417 ,           wr_2416 );
  not g1893( wr_2589 ,           wr_2588 );
  not g1894( wr_1686 ,           wr_1648 );
  not g1895( wr_2101 ,           wr_2065 );
  not g1896( wr_1538 ,           wr_1537 );
  not g1897( wr_1890 ,           wr_1853 );
  nor g1898( wr_1571 , wr_698  , wr_690  );
  nor g1899( wr_2490 , wr_265  , wr_243  );
  nor g1900( wr_2645 , wr_465  , wr_437  );
  nor g1901( wr_1556 , wr_1555 , wr_730  );
  nor g1902( wr_1614 , wr_1613 , wr_1602 );
  nor g1903( wr_2533 , wr_2532 , wr_2521 );
  nor g1904( wr_2688 , wr_2687 , wr_2676 );
  nor g1905( wr_1607 , wr_1606 , wr_1605 );
  nor g1906( wr_2526 , wr_2525 , wr_2524 );
  nor g1907( wr_2681 , wr_2680 , wr_2679 );
  not g1908( wr_1631 ,           wr_1630 );
  not g1909( wr_2550 ,           wr_2549 );
  not g1910( wr_2705 ,           wr_2704 );
  nor g1911( wr_1570 , wr_1569 , wr_1567 );
  nor g1912( wr_727  , wr_726  , wr_647  );
  not g1913( wr_2781 ,           wr_2780 );
  not g1914( wr_2959 ,           wr_2958 );
  not g1915( wr_3102 ,           wr_3101 );
  not g1916( wr_3279 ,           wr_3278 );
  nor g1917( wr_736  , wr_735  , wr_657  );
  not g1918( wr_2721 ,           wr_2720 );
  not g1919( wr_2908 ,           wr_2907 );
  not g1920( wr_3043 ,           wr_3042 );
  not g1921( wr_3228 ,           wr_3227 );
  nor g1922( wr_1521 , wr_1520 , wr_637  );
  nor g1923( wr_2361 , wr_2360 , wr_324  );
  nor g1924( wr_2423 , wr_2422 , wr_208  );
  nor g1925( wr_2595 , wr_2594 , wr_528  );
  nor g1926( wr_2768 , wr_2767 , wr_324  );
  nor g1927( wr_2946 , wr_2945 , wr_208  );
  nor g1928( wr_3089 , wr_3088 , wr_528  );
  nor g1929( wr_3266 , wr_3265 , wr_637  );
  nor g1930( wr_346  , wr_345  , wr_334  );
  nor g1931( wr_416  , wr_415  , wr_309  );
  nor g1932( wr_550  , wr_549  , wr_538  );
  nor g1933( wr_677  , wr_676  , wr_513  );
  nor g1934( wr_700  , wr_699  , wr_601  );
  not g1935( wr_1592 ,           wr_1591 );
  not g1936( wr_2511 ,           wr_2510 );
  not g1937( wr_2666 ,           wr_2665 );
  not g1938( wr_2825 ,           wr_2823 );
  not g1939( wr_3146 ,           wr_3144 );
  not g1940( wr_3323 ,           wr_3321 );
  nor g1941( wr_287  , wr_286  , wr_282  );
  nor g1942( wr_355  , wr_354  , wr_295  );
  nor g1943( wr_488  , wr_487  , wr_483  );
  nor g1944( wr_559  , wr_558  , wr_499  );
  nor g1945( wr_2824 , wr_2823 , wr_2545 );
  not g1946( wr_2852 ,           wr_2851 );
  nor g1947( wr_3145 , wr_3144 , wr_2700 );
  not g1948( wr_3173 ,           wr_3172 );
  nor g1949( wr_3322 , wr_3321 , wr_1626 );
  not g1950( wr_3350 ,           wr_3349 );
  nor g1951( wr_1447 , wr_1446 , wr_411  );
  nor g1952( wr_1484 , wr_1483 , wr_672  );
  nor g1953( wr_2857 , wr_2856 , wr_2855 );
  nor g1954( wr_3178 , wr_3177 , wr_3176 );
  nor g1955( wr_3355 , wr_3354 , wr_3353 );
  nor g1956( wr_267  , wr_266  , wr_239  );
  nor g1957( wr_467  , wr_466  , wr_431  );
  nor g1958( wr_616  , wr_615  , wr_581  );
  nor g1959( wr_662  , wr_661  , wr_627  );
  nor g1960( wr_1395 , wr_1394 , wr_1281 );
  not g1961( wr_2793 ,           wr_2777 );
  not g1962( wr_2971 ,           wr_2955 );
  not g1963( wr_3114 ,           wr_3098 );
  not g1964( wr_3291 ,           wr_3275 );
  nor g1965( wr_1438 , wr_1437 , wr_253  );
  nor g1966( wr_1457 , wr_1456 , wr_450  );
  nor g1967( wr_1404 , wr_1403 , wr_1312 );
  nor g1968( wr_1468 , wr_1467 , wr_611  );
  nor g1969( wr_1474 , wr_1473 , wr_162  );
  nor g1970( wr_387  , wr_386  , wr_215  );
  nor g1971( wr_972  , wr_971  , wr_958  );
  nor g1972( wr_1042 , wr_1041 , wr_1037 );
  nor g1973( wr_1345 , wr_1344 , wr_1340 );
  nor g1974( wr_1368 , wr_1367 , wr_1251 );
  nor g1975( wr_227  , wr_226  , wr_201  );
  nor g1976( wr_825  , wr_824  , wr_787  );
  nor g1977( wr_1194 , wr_1193 , wr_1180 );
  nor g1978( wr_1428 , wr_1427 , wr_194  );
  nor g1979( wr_396  , wr_395  , wr_222  );
  nor g1980( wr_901  , wr_900  , wr_863  );
  nor g1981( wr_981  , wr_980  , wr_913  );
  nor g1982( wr_1122 , wr_1121 , wr_1082 );
  nor g1983( wr_1771 , wr_1770 , wr_1766 );
  nor g1984( wr_1779 , wr_1778 , wr_1775 );
  nor g1985( wr_1822 , wr_1821 , wr_1817 );
  nor g1986( wr_1830 , wr_1829 , wr_1826 );
  nor g1987( wr_2184 , wr_2183 , wr_2179 );
  nor g1988( wr_2192 , wr_2191 , wr_2188 );
  nor g1989( wr_2233 , wr_2232 , wr_2228 );
  nor g1990( wr_2241 , wr_2240 , wr_2237 );
  nor g1991( wr_1203 , wr_1202 , wr_1135 );
  nor g1992( wr_881  , wr_880  , wr_841  );
  nor g1993( wr_1268 , wr_1267 , wr_1227 );
  nor g1994( wr_1329 , wr_1328 , wr_1288 );
  nor g1995( wr_1715 , wr_1714 , wr_1710 );
  nor g1996( wr_1723 , wr_1722 , wr_1719 );
  nor g1997( wr_1984 , wr_1983 , wr_1979 );
  nor g1998( wr_1992 , wr_1991 , wr_1988 );
  nor g1999( wr_2034 , wr_2033 , wr_2029 );
  nor g2000( wr_2042 , wr_2041 , wr_2038 );
  nor g2001( wr_2131 , wr_2130 , wr_2126 );
  nor g2002( wr_2139 , wr_2138 , wr_2135 );
  nor g2003( wr_1013 , wr_1012 , wr_778  );
  nor g2004( wr_1101 , wr_1100 , wr_1059 );
  nor g2005( wr_1673 , wr_1672 , wr_1668 );
  nor g2006( wr_1681 , wr_1680 , wr_1677 );
  nor g2007( wr_1929 , wr_1928 , wr_1924 );
  nor g2008( wr_1937 , wr_1936 , wr_1933 );
  nor g2009( wr_2088 , wr_2087 , wr_2083 );
  nor g2010( wr_2096 , wr_2095 , wr_2092 );
  nor g2011( wr_1022 , wr_1021 , wr_809  );
  nor g2012( wr_1516 , wr_1515 , wr_164  );
  nor g2013( wr_1877 , wr_1876 , wr_1872 );
  nor g2014( wr_1885 , wr_1884 , wr_1881 );
  nor g2015( wr_1539 , wr_1538 , wr_162  );
  not g2016( wr_1572 ,           wr_1571 );
  not g2017( wr_2491 ,           wr_2490 );
  not g2018( wr_2646 ,           wr_2645 );
  not g2019( wr_1557 ,           wr_1556 );
  not g2020( wr_1615 ,           wr_1614 );
  not g2021( wr_2534 ,           wr_2533 );
  not g2022( wr_2689 ,           wr_2688 );
  nor g2023( wr_1608 , wr_1607 , wr_1604 );
  nor g2024( wr_1617 , wr_1614 , wr_1605 );
  nor g2025( wr_2527 , wr_2526 , wr_2523 );
  nor g2026( wr_2536 , wr_2533 , wr_2524 );
  nor g2027( wr_2682 , wr_2681 , wr_2678 );
  nor g2028( wr_2691 , wr_2688 , wr_2679 );
  not g2029( G397    ,           wr_1570 );
  not g2030( wr_728  ,           wr_727  );
  nor g2031( wr_2782 , wr_2781 , wr_315  );
  nor g2032( wr_2960 , wr_2959 , wr_376  );
  nor g2033( wr_3103 , wr_3102 , wr_519  );
  nor g2034( wr_3280 , wr_3279 , wr_716  );
  nor g2035( wr_2722 , wr_2721 , wr_2374 );
  nor g2036( wr_2909 , wr_2908 , wr_2436 );
  nor g2037( wr_3044 , wr_3043 , wr_2608 );
  nor g2038( wr_3229 , wr_3228 , wr_1534 );
  nor g2039( wr_2769 , wr_2768 , wr_2361 );
  nor g2040( wr_2947 , wr_2946 , wr_2423 );
  nor g2041( wr_3090 , wr_3089 , wr_2595 );
  nor g2042( wr_3267 , wr_3266 , wr_1521 );
  not g2043( wr_347  ,           wr_346  );
  not g2044( wr_417  ,           wr_416  );
  not g2045( wr_551  ,           wr_550  );
  not g2046( wr_678  ,           wr_677  );
  nor g2047( wr_706  , wr_705  , wr_700  );
  nor g2048( wr_1593 , wr_1592 , wr_690  );
  nor g2049( wr_2512 , wr_2511 , wr_243  );
  nor g2050( wr_2667 , wr_2666 , wr_437  );
  nor g2051( wr_2712 , wr_2361 , wr_2351 );
  nor g2052( wr_2899 , wr_2423 , wr_2413 );
  nor g2053( wr_3034 , wr_2595 , wr_2585 );
  nor g2054( wr_3219 , wr_1521 , wr_1511 );
  nor g2055( wr_2826 , wr_2825 , wr_2547 );
  nor g2056( wr_3147 , wr_3146 , wr_2702 );
  nor g2057( wr_3324 , wr_3323 , wr_1628 );
  not g2058( wr_288  ,           wr_287  );
  not g2059( wr_489  ,           wr_488  );
  nor g2060( wr_2853 , wr_2852 , wr_270  );
  nor g2061( wr_3174 , wr_3173 , wr_470  );
  nor g2062( wr_3351 , wr_3350 , wr_703  );
  not g2063( wr_1448 ,           wr_1447 );
  not g2064( wr_1485 ,           wr_1484 );
  not g2065( wr_2858 ,           wr_2857 );
  not g2066( wr_3179 ,           wr_3178 );
  not g2067( wr_3356 ,           wr_3355 );
  nor g2068( wr_273  , wr_272  , wr_267  );
  nor g2069( wr_473  , wr_472  , wr_467  );
  not g2070( wr_617  ,           wr_616  );
  not g2071( wr_663  ,           wr_662  );
  not g2072( wr_1396 ,           wr_1395 );
  not g2073( wr_1439 ,           wr_1438 );
  not g2074( wr_1458 ,           wr_1457 );
  not g2075( wr_1469 ,           wr_1468 );
  not g2076( wr_1475 ,           wr_1474 );
  not g2077( wr_388  ,           wr_387  );
  not g2078( wr_973  ,           wr_972  );
  not g2079( wr_1043 ,           wr_1042 );
  not g2080( wr_1346 ,           wr_1345 );
  nor g2081( wr_1374 , wr_1373 , wr_1368 );
  not g2082( wr_228  ,           wr_227  );
  not g2083( wr_826  ,           wr_825  );
  not g2084( wr_1195 ,           wr_1194 );
  not g2085( wr_1429 ,           wr_1428 );
  not g2086( wr_902  ,           wr_901  );
  not g2087( wr_1123 ,           wr_1122 );
  not g2088( wr_1772 ,           wr_1771 );
  not g2089( wr_1780 ,           wr_1779 );
  not g2090( wr_1823 ,           wr_1822 );
  not g2091( wr_1831 ,           wr_1830 );
  not g2092( wr_2185 ,           wr_2184 );
  not g2093( wr_2193 ,           wr_2192 );
  not g2094( wr_2234 ,           wr_2233 );
  not g2095( wr_2242 ,           wr_2241 );
  nor g2096( wr_887  , wr_886  , wr_881  );
  not g2097( wr_1269 ,           wr_1268 );
  not g2098( wr_1330 ,           wr_1329 );
  not g2099( wr_1716 ,           wr_1715 );
  not g2100( wr_1724 ,           wr_1723 );
  not g2101( wr_1985 ,           wr_1984 );
  not g2102( wr_1993 ,           wr_1992 );
  not g2103( wr_2035 ,           wr_2034 );
  not g2104( wr_2043 ,           wr_2042 );
  not g2105( wr_2132 ,           wr_2131 );
  not g2106( wr_2140 ,           wr_2139 );
  not g2107( wr_1014 ,           wr_1013 );
  nor g2108( wr_1107 , wr_1106 , wr_1101 );
  not g2109( wr_1674 ,           wr_1673 );
  not g2110( wr_1682 ,           wr_1681 );
  not g2111( wr_1930 ,           wr_1929 );
  not g2112( wr_1938 ,           wr_1937 );
  not g2113( wr_2089 ,           wr_2088 );
  not g2114( wr_2097 ,           wr_2096 );
  not g2115( wr_1517 ,           wr_1516 );
  not g2116( wr_1878 ,           wr_1877 );
  not g2117( wr_1886 ,           wr_1885 );
  nor g2118( wr_1543 , wr_1542 , wr_1539 );
  nor g2119( wr_1573 , wr_1572 , wr_703  );
  nor g2120( wr_2492 , wr_2491 , wr_270  );
  nor g2121( wr_2647 , wr_2646 , wr_470  );
  nor g2122( wr_1558 , wr_1557 , wr_1540 );
  nor g2123( wr_1616 , wr_1615 , wr_591  );
  nor g2124( wr_2535 , wr_2534 , wr_257  );
  nor g2125( wr_2690 , wr_2689 , wr_455  );
  not g2126( wr_1609 ,           wr_1608 );
  not g2127( wr_2528 ,           wr_2527 );
  not g2128( wr_2683 ,           wr_2682 );
  nor g2129( wr_729  , wr_728  , wr_637  );
  not g2130( wr_2783 ,           wr_2782 );
  not g2131( wr_2961 ,           wr_2960 );
  not g2132( wr_3104 ,           wr_3103 );
  not g2133( wr_3281 ,           wr_3280 );
  not g2134( wr_2723 ,           wr_2722 );
  not g2135( wr_2910 ,           wr_2909 );
  not g2136( wr_3045 ,           wr_3044 );
  not g2137( wr_3230 ,           wr_3229 );
  nor g2138( wr_2725 , wr_2722 , wr_341  );
  not g2139( wr_2770 ,           wr_2769 );
  nor g2140( wr_2912 , wr_2909 , wr_382  );
  not g2141( wr_2948 ,           wr_2947 );
  nor g2142( wr_3047 , wr_3044 , wr_545  );
  not g2143( wr_3091 ,           wr_3090 );
  nor g2144( wr_3232 , wr_3229 , wr_722  );
  not g2145( wr_3268 ,           wr_3267 );
  nor g2146( wr_348  , wr_347  , wr_324  );
  nor g2147( wr_418  , wr_417  , wr_411  );
  nor g2148( wr_552  , wr_551  , wr_528  );
  nor g2149( wr_679  , wr_678  , wr_672  );
  not g2150( wr_707  ,           wr_706  );
  not g2151( wr_1594 ,           wr_1593 );
  not g2152( wr_2513 ,           wr_2512 );
  not g2153( wr_2668 ,           wr_2667 );
  not g2154( wr_2713 ,           wr_2712 );
  not g2155( wr_2900 ,           wr_2899 );
  not g2156( wr_3035 ,           wr_3034 );
  not g2157( wr_3220 ,           wr_3219 );
  nor g2158( wr_2827 , wr_2826 , wr_2824 );
  nor g2159( wr_3148 , wr_3147 , wr_3145 );
  nor g2160( wr_3325 , wr_3324 , wr_3322 );
  not g2161( wr_2854 ,           wr_2853 );
  not g2162( wr_3175 ,           wr_3174 );
  not g2163( wr_3352 ,           wr_3351 );
  nor g2164( wr_1449 , wr_1448 , wr_334  );
  nor g2165( wr_1486 , wr_1485 , wr_538  );
  nor g2166( wr_2860 , wr_2857 , wr_2853 );
  nor g2167( wr_3181 , wr_3178 , wr_3174 );
  nor g2168( wr_3358 , wr_3355 , wr_3351 );
  not g2169( wr_274  ,           wr_273  );
  not g2170( wr_474  ,           wr_473  );
  nor g2171( wr_664  , wr_663  , wr_162  );
  nor g2172( wr_1397 , wr_1396 , wr_1300 );
  nor g2173( wr_1476 , wr_1475 , wr_647  );
  nor g2174( wr_389  , wr_388  , wr_208  );
  nor g2175( wr_974  , wr_973  , wr_946  );
  nor g2176( wr_1044 , wr_1043 , wr_958  );
  nor g2177( wr_1347 , wr_1346 , wr_1180 );
  not g2178( wr_1375 ,           wr_1374 );
  nor g2179( wr_229  , wr_228  , wr_194  );
  nor g2180( wr_827  , wr_826  , wr_778  );
  nor g2181( wr_1196 , wr_1195 , wr_1168 );
  nor g2182( wr_1430 , wr_1429 , wr_215  );
  nor g2183( wr_1781 , wr_1780 , wr_1772 );
  nor g2184( wr_1832 , wr_1831 , wr_1823 );
  nor g2185( wr_2194 , wr_2193 , wr_2185 );
  nor g2186( wr_2243 , wr_2242 , wr_2234 );
  not g2187( wr_888  ,           wr_887  );
  nor g2188( wr_1331 , wr_1330 , wr_1281 );
  nor g2189( wr_1725 , wr_1724 , wr_1716 );
  nor g2190( wr_1994 , wr_1993 , wr_1985 );
  nor g2191( wr_2044 , wr_2043 , wr_2035 );
  nor g2192( wr_2141 , wr_2140 , wr_2132 );
  nor g2193( wr_1015 , wr_1014 , wr_798  );
  not g2194( wr_1108 ,           wr_1107 );
  nor g2195( wr_1683 , wr_1682 , wr_1674 );
  nor g2196( wr_1939 , wr_1938 , wr_1930 );
  nor g2197( wr_2098 , wr_2097 , wr_2089 );
  nor g2198( wr_1518 , wr_1517 , wr_162  );
  nor g2199( wr_1887 , wr_1886 , wr_1878 );
  not g2200( wr_1544 ,           wr_1543 );
  not g2201( wr_1576 ,           wr_1573 );
  not g2202( wr_2495 ,           wr_2492 );
  not g2203( wr_2650 ,           wr_2647 );
  nor g2204( wr_1574 , wr_1573 , wr_601  );
  nor g2205( wr_2493 , wr_2492 , wr_239  );
  nor g2206( wr_2648 , wr_2647 , wr_431  );
  not g2207( wr_1559 ,           wr_1558 );
  nor g2208( wr_1618 , wr_1617 , wr_1616 );
  nor g2209( wr_2537 , wr_2536 , wr_2535 );
  nor g2210( wr_2692 , wr_2691 , wr_2690 );
  nor g2211( wr_1562 , wr_1558 , wr_1561 );
  nor g2212( wr_737  , wr_736  , wr_729  );
  nor g2213( wr_2784 , wr_2783 , wr_2374 );
  nor g2214( wr_2962 , wr_2961 , wr_2436 );
  nor g2215( wr_3105 , wr_3104 , wr_2608 );
  nor g2216( wr_3282 , wr_3281 , wr_1534 );
  nor g2217( wr_2724 , wr_2723 , wr_340  );
  nor g2218( wr_2911 , wr_2910 , wr_381  );
  nor g2219( wr_3046 , wr_3045 , wr_544  );
  nor g2220( wr_3231 , wr_3230 , wr_721  );
  nor g2221( wr_2771 , wr_2770 , wr_2351 );
  nor g2222( wr_2949 , wr_2948 , wr_2413 );
  nor g2223( wr_3092 , wr_3091 , wr_2585 );
  nor g2224( wr_3269 , wr_3268 , wr_1511 );
  nor g2225( wr_356  , wr_355  , wr_348  );
  not g2226( wr_419  ,           wr_418  );
  nor g2227( wr_560  , wr_559  , wr_552  );
  not g2228( wr_680  ,           wr_679  );
  nor g2229( wr_708  , wr_707  , wr_693  );
  nor g2230( wr_1595 , wr_1594 , wr_703  );
  nor g2231( wr_2514 , wr_2513 , wr_270  );
  nor g2232( wr_2669 , wr_2668 , wr_470  );
  nor g2233( wr_2714 , wr_2713 , wr_301  );
  nor g2234( wr_2901 , wr_2900 , wr_372  );
  nor g2235( wr_3036 , wr_3035 , wr_505  );
  nor g2236( wr_3221 , wr_3220 , wr_712  );
  not g2237( wr_2828 ,           wr_2827 );
  not g2238( wr_3149 ,           wr_3148 );
  not g2239( wr_3326 ,           wr_3325 );
  nor g2240( wr_2859 , wr_2858 , wr_2854 );
  nor g2241( wr_3180 , wr_3179 , wr_3175 );
  nor g2242( wr_3357 , wr_3356 , wr_3352 );
  not g2243( wr_1450 ,           wr_1449 );
  not g2244( wr_1487 ,           wr_1486 );
  nor g2245( wr_275  , wr_274  , wr_246  );
  nor g2246( wr_475  , wr_474  , wr_440  );
  not g2247( wr_665  ,           wr_664  );
  nor g2248( wr_1405 , wr_1404 , wr_1397 );
  not g2249( wr_1477 ,           wr_1476 );
  nor g2250( wr_397  , wr_396  , wr_389  );
  nor g2251( wr_982  , wr_981  , wr_974  );
  not g2252( wr_1045 ,           wr_1044 );
  not g2253( wr_1348 ,           wr_1347 );
  nor g2254( wr_1376 , wr_1375 , wr_1361 );
  not g2255( wr_230  ,           wr_229  );
  not g2256( wr_828  ,           wr_827  );
  nor g2257( wr_1204 , wr_1203 , wr_1196 );
  not g2258( wr_1431 ,           wr_1430 );
  not g2259( wr_1782 ,           wr_1781 );
  not g2260( wr_1833 ,           wr_1832 );
  not g2261( wr_2195 ,           wr_2194 );
  not g2262( wr_2244 ,           wr_2243 );
  nor g2263( wr_1785 , wr_1781 , wr_1784 );
  nor g2264( wr_1836 , wr_1832 , wr_1835 );
  nor g2265( wr_2198 , wr_2194 , wr_2197 );
  nor g2266( wr_2247 , wr_2243 , wr_2246 );
  nor g2267( wr_889  , wr_888  , wr_852  );
  not g2268( wr_1332 ,           wr_1331 );
  not g2269( wr_1726 ,           wr_1725 );
  not g2270( wr_1995 ,           wr_1994 );
  not g2271( wr_2045 ,           wr_2044 );
  not g2272( wr_2142 ,           wr_2141 );
  nor g2273( wr_1023 , wr_1022 , wr_1015 );
  nor g2274( wr_1109 , wr_1108 , wr_1070 );
  nor g2275( wr_1729 , wr_1725 , wr_1728 );
  nor g2276( wr_1998 , wr_1994 , wr_1997 );
  nor g2277( wr_2048 , wr_2044 , wr_2047 );
  nor g2278( wr_2145 , wr_2141 , wr_2144 );
  not g2279( wr_1684 ,           wr_1683 );
  not g2280( wr_1940 ,           wr_1939 );
  not g2281( wr_2099 ,           wr_2098 );
  nor g2282( wr_1687 , wr_1683 , wr_1686 );
  nor g2283( wr_1943 , wr_1939 , wr_1942 );
  nor g2284( wr_2102 , wr_2098 , wr_2101 );
  nor g2285( wr_1522 , wr_1521 , wr_1518 );
  not g2286( wr_1888 ,           wr_1887 );
  nor g2287( wr_1891 , wr_1887 , wr_1890 );
  nor g2288( wr_1545 , wr_1544 , wr_716  );
  nor g2289( wr_1577 , wr_1576 , wr_1575 );
  nor g2290( wr_2496 , wr_2495 , wr_2494 );
  nor g2291( wr_2651 , wr_2650 , wr_2649 );
  nor g2292( wr_1560 , wr_1559 , wr_637  );
  not g2293( wr_738  ,           wr_737  );
  not g2294( wr_2787 ,           wr_2784 );
  not g2295( wr_2965 ,           wr_2962 );
  not g2296( wr_3108 ,           wr_3105 );
  not g2297( wr_3285 ,           wr_3282 );
  nor g2298( wr_2726 , wr_2725 , wr_2724 );
  nor g2299( wr_2786 , wr_2785 , wr_2784 );
  nor g2300( wr_2913 , wr_2912 , wr_2911 );
  nor g2301( wr_2964 , wr_2963 , wr_2962 );
  nor g2302( wr_3048 , wr_3047 , wr_3046 );
  nor g2303( wr_3107 , wr_3106 , wr_3105 );
  nor g2304( wr_3233 , wr_3232 , wr_3231 );
  nor g2305( wr_3284 , wr_3283 , wr_3282 );
  not g2306( wr_2772 ,           wr_2771 );
  not g2307( wr_2950 ,           wr_2949 );
  not g2308( wr_3093 ,           wr_3092 );
  not g2309( wr_3270 ,           wr_3269 );
  not g2310( wr_357  ,           wr_356  );
  nor g2311( wr_420  , wr_419  , wr_288  );
  not g2312( wr_561  ,           wr_560  );
  nor g2313( wr_681  , wr_680  , wr_489  );
  not g2314( wr_709  ,           wr_708  );
  not g2315( wr_1596 ,           wr_1595 );
  not g2316( wr_2515 ,           wr_2514 );
  not g2317( wr_2670 ,           wr_2669 );
  not g2318( wr_2715 ,           wr_2714 );
  not g2319( wr_2902 ,           wr_2901 );
  not g2320( wr_3037 ,           wr_3036 );
  not g2321( wr_3222 ,           wr_3221 );
  nor g2322( wr_2829 , wr_2828 , wr_2514 );
  nor g2323( wr_3150 , wr_3149 , wr_2669 );
  nor g2324( wr_3327 , wr_3326 , wr_1595 );
  nor g2325( wr_2861 , wr_2860 , wr_2859 );
  nor g2326( wr_3182 , wr_3181 , wr_3180 );
  nor g2327( wr_3359 , wr_3358 , wr_3357 );
  nor g2328( wr_1451 , wr_1450 , wr_1439 );
  nor g2329( wr_1488 , wr_1487 , wr_1458 );
  not g2330( wr_276  ,           wr_275  );
  not g2331( wr_476  ,           wr_475  );
  nor g2332( wr_666  , wr_665  , wr_617  );
  not g2333( wr_1406 ,           wr_1405 );
  nor g2334( wr_1478 , wr_1477 , wr_1469 );
  nor g2335( wr_1581 , wr_665  , wr_164  );
  not g2336( wr_398  ,           wr_397  );
  not g2337( wr_983  ,           wr_982  );
  nor g2338( wr_1046 , wr_1045 , wr_902  );
  nor g2339( wr_1349 , wr_1348 , wr_1123 );
  not g2340( wr_1377 ,           wr_1376 );
  nor g2341( wr_231  , wr_230  , wr_183  );
  nor g2342( wr_829  , wr_828  , wr_767  );
  not g2343( wr_1205 ,           wr_1204 );
  nor g2344( wr_1432 , wr_1431 , wr_183  );
  nor g2345( wr_1783 , wr_1782 , wr_1741 );
  nor g2346( wr_1834 , wr_1833 , wr_1797 );
  nor g2347( wr_2196 , wr_2195 , wr_2157 );
  nor g2348( wr_2245 , wr_2244 , wr_2210 );
  nor g2349( wr_3079 , wr_1477 , wr_164  );
  not g2350( wr_890  ,           wr_889  );
  nor g2351( wr_1333 , wr_1332 , wr_1269 );
  nor g2352( wr_1727 , wr_1726 , wr_1697 );
  nor g2353( wr_1996 , wr_1995 , wr_1955 );
  nor g2354( wr_2046 , wr_2045 , wr_2010 );
  nor g2355( wr_2143 , wr_2142 , wr_2112 );
  not g2356( wr_1024 ,           wr_1023 );
  not g2357( wr_1110 ,           wr_1109 );
  nor g2358( wr_1685 , wr_1684 , wr_1648 );
  nor g2359( wr_1941 , wr_1940 , wr_1905 );
  nor g2360( wr_2100 , wr_2099 , wr_2065 );
  nor g2361( wr_2314 , wr_1332 , wr_1335 );
  not g2362( wr_1523 ,           wr_1522 );
  nor g2363( wr_1889 , wr_1888 , wr_1853 );
  not g2364( wr_1546 ,           wr_1545 );
  nor g2365( wr_1578 , wr_1577 , wr_1574 );
  nor g2366( wr_1598 , wr_1595 , wr_1575 );
  nor g2367( wr_2497 , wr_2496 , wr_2493 );
  nor g2368( wr_2517 , wr_2514 , wr_2494 );
  nor g2369( wr_2652 , wr_2651 , wr_2648 );
  nor g2370( wr_2672 , wr_2669 , wr_2649 );
  nor g2371( wr_1563 , wr_1562 , wr_1560 );
  nor g2372( wr_739  , wr_738  , wr_720  );
  nor g2373( wr_2789 , wr_2788 , wr_2787 );
  nor g2374( wr_2967 , wr_2966 , wr_2965 );
  nor g2375( wr_3110 , wr_3109 , wr_3108 );
  nor g2376( wr_3287 , wr_3286 , wr_3285 );
  not g2377( wr_2727 ,           wr_2726 );
  not g2378( wr_2914 ,           wr_2913 );
  not g2379( wr_3049 ,           wr_3048 );
  not g2380( wr_3234 ,           wr_3233 );
  nor g2381( wr_2729 , wr_2726 , wr_2718 );
  nor g2382( wr_2773 , wr_2772 , wr_301  );
  nor g2383( wr_2916 , wr_2913 , wr_2905 );
  nor g2384( wr_2951 , wr_2950 , wr_372  );
  nor g2385( wr_3051 , wr_3048 , wr_3040 );
  nor g2386( wr_3094 , wr_3093 , wr_505  );
  nor g2387( wr_3236 , wr_3233 , wr_3225 );
  nor g2388( wr_3271 , wr_3270 , wr_712  );
  nor g2389( wr_358  , wr_357  , wr_319  );
  not g2390( wr_421  ,           wr_420  );
  nor g2391( wr_562  , wr_561  , wr_523  );
  not g2392( wr_682  ,           wr_681  );
  nor g2393( wr_710  , wr_709  , wr_692  );
  nor g2394( wr_2716 , wr_2715 , wr_317  );
  nor g2395( wr_2830 , wr_2827 , wr_2515 );
  nor g2396( wr_2903 , wr_2902 , wr_378  );
  nor g2397( wr_3038 , wr_3037 , wr_521  );
  nor g2398( wr_3151 , wr_3148 , wr_2670 );
  nor g2399( wr_3223 , wr_3222 , wr_718  );
  nor g2400( wr_3328 , wr_3325 , wr_1596 );
  not g2401( wr_2862 ,           wr_2861 );
  not g2402( wr_3183 ,           wr_3182 );
  not g2403( wr_3360 ,           wr_3359 );
  not g2404( wr_1452 ,           wr_1451 );
  not g2405( wr_1489 ,           wr_1488 );
  nor g2406( wr_2864 , wr_2861 , wr_2554 );
  nor g2407( wr_3185 , wr_3182 , wr_2709 );
  nor g2408( wr_3362 , wr_3359 , wr_1635 );
  nor g2409( wr_277  , wr_276  , wr_245  );
  nor g2410( wr_477  , wr_476  , wr_439  );
  not g2411( wr_667  ,           wr_666  );
  nor g2412( wr_1407 , wr_1406 , wr_1388 );
  not g2413( wr_1479 ,           wr_1478 );
  nor g2414( wr_399  , wr_398  , wr_380  );
  nor g2415( wr_984  , wr_983  , wr_941  );
  not g2416( wr_1047 ,           wr_1046 );
  not g2417( wr_1350 ,           wr_1349 );
  nor g2418( wr_1378 , wr_1377 , wr_1360 );
  not g2419( wr_232  ,           wr_231  );
  not g2420( wr_830  ,           wr_829  );
  nor g2421( wr_1206 , wr_1205 , wr_1163 );
  not g2422( wr_1433 ,           wr_1432 );
  nor g2423( wr_1786 , wr_1785 , wr_1783 );
  nor g2424( wr_1837 , wr_1836 , wr_1834 );
  nor g2425( wr_2199 , wr_2198 , wr_2196 );
  nor g2426( wr_2248 , wr_2247 , wr_2245 );
  nor g2427( wr_891  , wr_890  , wr_851  );
  not g2428( wr_1334 ,           wr_1333 );
  nor g2429( wr_1730 , wr_1729 , wr_1727 );
  nor g2430( wr_1999 , wr_1998 , wr_1996 );
  nor g2431( wr_2049 , wr_2048 , wr_2046 );
  nor g2432( wr_2146 , wr_2145 , wr_2143 );
  nor g2433( wr_1025 , wr_1024 , wr_1006 );
  nor g2434( wr_1111 , wr_1110 , wr_1069 );
  nor g2435( wr_1688 , wr_1687 , wr_1685 );
  nor g2436( wr_1944 , wr_1943 , wr_1941 );
  nor g2437( wr_2103 , wr_2102 , wr_2100 );
  nor g2438( wr_1524 , wr_1523 , wr_1511 );
  nor g2439( wr_1892 , wr_1891 , wr_1889 );
  nor g2440( wr_1547 , wr_1546 , wr_1534 );
  nor g2441( wr_1597 , wr_1596 , wr_601  );
  nor g2442( wr_2516 , wr_2515 , wr_239  );
  nor g2443( wr_2671 , wr_2670 , wr_431  );
  not g2444( wr_1579 ,           wr_1578 );
  not g2445( wr_2498 ,           wr_2497 );
  not g2446( wr_2653 ,           wr_2652 );
  not g2447( G394    ,           wr_1563 );
  not g2448( wr_740  ,           wr_739  );
  nor g2449( wr_2790 , wr_2789 , wr_2786 );
  nor g2450( wr_2968 , wr_2967 , wr_2964 );
  nor g2451( wr_3111 , wr_3110 , wr_3107 );
  nor g2452( wr_3288 , wr_3287 , wr_3284 );
  nor g2453( wr_2728 , wr_2727 , wr_2719 );
  nor g2454( wr_2915 , wr_2914 , wr_2906 );
  nor g2455( wr_3050 , wr_3049 , wr_3041 );
  nor g2456( wr_3235 , wr_3234 , wr_3226 );
  not g2457( wr_2774 ,           wr_2773 );
  not g2458( wr_2952 ,           wr_2951 );
  not g2459( wr_3095 ,           wr_3094 );
  not g2460( wr_3272 ,           wr_3271 );
  not g2461( wr_359  ,           wr_358  );
  not g2462( wr_563  ,           wr_562  );
  not g2463( wr_711  ,           wr_710  );
  nor g2464( wr_2292 , wr_682  , wr_421  );
  not g2465( wr_2717 ,           wr_2716 );
  nor g2466( wr_2831 , wr_2830 , wr_2829 );
  not g2467( wr_2904 ,           wr_2903 );
  not g2468( wr_3039 ,           wr_3038 );
  nor g2469( wr_3152 , wr_3151 , wr_3150 );
  not g2470( wr_3224 ,           wr_3223 );
  nor g2471( wr_3329 , wr_3328 , wr_3327 );
  nor g2472( wr_2863 , wr_2862 , wr_282  );
  nor g2473( wr_3184 , wr_3183 , wr_483  );
  nor g2474( wr_3361 , wr_3360 , wr_581  );
  nor g2475( wr_2330 , wr_1489 , wr_1452 );
  not g2476( wr_278  ,           wr_277  );
  not g2477( wr_478  ,           wr_477  );
  not g2478( wr_1408 ,           wr_1407 );
  nor g2479( wr_2279 , wr_682  , wr_164  );
  nor g2480( wr_2758 , wr_1489 , wr_164  );
  not g2481( wr_400  ,           wr_399  );
  not g2482( wr_985  ,           wr_984  );
  not g2483( wr_1379 ,           wr_1378 );
  nor g2484( wr_2258 , wr_1350 , wr_1047 );
  nor g2485( wr_683  , wr_421  , wr_232  );
  not g2486( wr_1207 ,           wr_1206 );
  nor g2487( wr_1351 , wr_1047 , wr_830  );
  nor g2488( wr_1490 , wr_1452 , wr_1433 );
  nor g2489( wr_1838 , wr_1837 , wr_1786 );
  nor g2490( wr_2249 , wr_2248 , wr_2199 );
  not g2491( wr_892  ,           wr_891  );
  nor g2492( wr_2050 , wr_2049 , wr_1999 );
  not g2493( wr_1026 ,           wr_1025 );
  not g2494( wr_1112 ,           wr_1111 );
  not g2495( wr_1525 ,           wr_1524 );
  not g2496( wr_1548 ,           wr_1547 );
  nor g2497( wr_1599 , wr_1598 , wr_1597 );
  nor g2498( wr_2518 , wr_2517 , wr_2516 );
  nor g2499( wr_2673 , wr_2672 , wr_2671 );
  nor g2500( wr_1551 , wr_1547 , wr_1550 );
  nor g2501( wr_741  , wr_740  , wr_715  );
  not g2502( wr_2791 ,           wr_2790 );
  not g2503( wr_2969 ,           wr_2968 );
  not g2504( wr_3112 ,           wr_3111 );
  not g2505( wr_3289 ,           wr_3288 );
  nor g2506( wr_2730 , wr_2729 , wr_2728 );
  nor g2507( wr_2794 , wr_2790 , wr_2793 );
  nor g2508( wr_2917 , wr_2916 , wr_2915 );
  nor g2509( wr_2972 , wr_2968 , wr_2971 );
  nor g2510( wr_3052 , wr_3051 , wr_3050 );
  nor g2511( wr_3115 , wr_3111 , wr_3114 );
  nor g2512( wr_3237 , wr_3236 , wr_3235 );
  nor g2513( wr_3292 , wr_3288 , wr_3291 );
  nor g2514( wr_2775 , wr_2774 , wr_317  );
  nor g2515( wr_2953 , wr_2952 , wr_378  );
  nor g2516( wr_3096 , wr_3095 , wr_521  );
  nor g2517( wr_3273 , wr_3272 , wr_718  );
  nor g2518( wr_360  , wr_359  , wr_304  );
  nor g2519( wr_564  , wr_563  , wr_508  );
  not g2520( wr_2293 ,           wr_2292 );
  not g2521( wr_2832 ,           wr_2831 );
  not g2522( wr_3153 ,           wr_3152 );
  not g2523( wr_3330 ,           wr_3329 );
  nor g2524( wr_2834 , wr_2831 , wr_2554 );
  nor g2525( wr_3155 , wr_3152 , wr_2709 );
  nor g2526( wr_3332 , wr_3329 , wr_1635 );
  nor g2527( wr_2865 , wr_2864 , wr_2863 );
  nor g2528( wr_3186 , wr_3185 , wr_3184 );
  nor g2529( wr_3363 , wr_3362 , wr_3361 );
  not g2530( wr_2331 ,           wr_2330 );
  nor g2531( wr_1409 , wr_1408 , wr_1383 );
  not g2532( wr_2280 ,           wr_2279 );
  nor g2533( wr_2558 , wr_711  , wr_616  );
  not g2534( wr_2759 ,           wr_2758 );
  nor g2535( wr_401  , wr_400  , wr_375  );
  nor g2536( wr_986  , wr_985  , wr_924  );
  not g2537( wr_2259 ,           wr_2258 );
  not g2538( wr_684  ,           wr_683  );
  nor g2539( wr_1208 , wr_1207 , wr_1146 );
  not g2540( wr_1352 ,           wr_1351 );
  not g2541( wr_1491 ,           wr_1490 );
  nor g2542( wr_3078 , wr_1468 , wr_711  );
  not g2543( wr_1839 ,           wr_1838 );
  not g2544( wr_2250 ,           wr_2249 );
  not g2545( wr_2051 ,           wr_2050 );
  nor g2546( wr_1027 , wr_1026 , wr_1001 );
  nor g2547( wr_2312 , wr_1379 , wr_1268 );
  nor g2548( wr_1526 , wr_1525 , wr_712  );
  nor g2549( wr_2310 , wr_1122 , wr_1112 );
  nor g2550( wr_1549 , wr_1548 , wr_627  );
  not g2551( wr_742  ,           wr_741  );
  nor g2552( wr_2792 , wr_2791 , wr_2777 );
  nor g2553( wr_2970 , wr_2969 , wr_2955 );
  nor g2554( wr_3113 , wr_3112 , wr_3098 );
  nor g2555( wr_3290 , wr_3289 , wr_3275 );
  not g2556( wr_2731 ,           wr_2730 );
  not g2557( wr_2918 ,           wr_2917 );
  not g2558( wr_3053 ,           wr_3052 );
  not g2559( wr_3238 ,           wr_3237 );
  nor g2560( wr_2733 , wr_2730 , wr_2716 );
  not g2561( wr_2798 ,           wr_2775 );
  nor g2562( wr_2920 , wr_2917 , wr_2903 );
  not g2563( wr_2976 ,           wr_2953 );
  nor g2564( wr_3055 , wr_3052 , wr_3038 );
  not g2565( wr_3119 ,           wr_3096 );
  nor g2566( wr_3240 , wr_3237 , wr_3223 );
  not g2567( wr_3296 ,           wr_3273 );
  not g2568( wr_361  ,           wr_360  );
  not g2569( wr_565  ,           wr_564  );
  nor g2570( wr_2294 , wr_2293 , wr_164  );
  nor g2571( wr_2833 , wr_2832 , wr_282  );
  nor g2572( wr_3154 , wr_3153 , wr_483  );
  nor g2573( wr_3331 , wr_3330 , wr_581  );
  not g2574( wr_2866 ,           wr_2865 );
  not g2575( wr_3187 ,           wr_3186 );
  not g2576( wr_3364 ,           wr_3363 );
  nor g2577( wr_2332 , wr_2331 , wr_164  );
  nor g2578( wr_2868 , wr_2865 , wr_2541 );
  nor g2579( wr_3189 , wr_3186 , wr_2696 );
  nor g2580( wr_3366 , wr_3363 , wr_1622 );
  not g2581( wr_1410 ,           wr_1409 );
  nor g2582( wr_2281 , wr_2280 , wr_667  );
  nor g2583( wr_2760 , wr_2759 , wr_1479 );
  not g2584( wr_402  ,           wr_401  );
  not g2585( wr_987  ,           wr_986  );
  nor g2586( wr_2260 , wr_2259 , wr_1335 );
  nor g2587( wr_685  , wr_684  , wr_682  );
  not g2588( wr_1209 ,           wr_1208 );
  nor g2589( wr_1353 , wr_1352 , wr_1350 );
  nor g2590( wr_1492 , wr_1491 , wr_1489 );
  nor g2591( wr_1840 , wr_1839 , wr_1730 );
  nor g2592( wr_2251 , wr_2250 , wr_2146 );
  nor g2593( wr_2052 , wr_2051 , wr_1944 );
  not g2594( wr_1028 ,           wr_1027 );
  not g2595( wr_1527 ,           wr_1526 );
  nor g2596( wr_1552 , wr_1551 , wr_1549 );
  nor g2597( wr_743  , wr_742  , wr_714  );
  nor g2598( wr_2795 , wr_2794 , wr_2792 );
  nor g2599( wr_2973 , wr_2972 , wr_2970 );
  nor g2600( wr_3116 , wr_3115 , wr_3113 );
  nor g2601( wr_3293 , wr_3292 , wr_3290 );
  nor g2602( wr_2732 , wr_2731 , wr_2717 );
  nor g2603( wr_2919 , wr_2918 , wr_2904 );
  nor g2604( wr_3054 , wr_3053 , wr_3039 );
  nor g2605( wr_3239 , wr_3238 , wr_3224 );
  nor g2606( wr_362  , wr_361  , wr_303  );
  nor g2607( wr_566  , wr_565  , wr_507  );
  not g2608( wr_2295 ,           wr_2294 );
  nor g2609( wr_2835 , wr_2834 , wr_2833 );
  nor g2610( wr_3156 , wr_3155 , wr_3154 );
  nor g2611( wr_3333 , wr_3332 , wr_3331 );
  nor g2612( wr_2867 , wr_2866 , wr_253  );
  nor g2613( wr_3188 , wr_3187 , wr_450  );
  nor g2614( wr_3365 , wr_3364 , wr_611  );
  not g2615( wr_2333 ,           wr_2332 );
  nor g2616( wr_1411 , wr_1410 , wr_1382 );
  nor g2617( wr_403  , wr_402  , wr_374  );
  nor g2618( wr_988  , wr_987  , wr_923  );
  not g2619( wr_2261 ,           wr_2260 );
  not g2620( wr_686  ,           wr_685  );
  nor g2621( wr_1210 , wr_1209 , wr_1145 );
  not g2622( wr_1354 ,           wr_1353 );
  not g2623( wr_1493 ,           wr_1492 );
  not g2624( wr_1841 ,           wr_1840 );
  not g2625( wr_2252 ,           wr_2251 );
  not g2626( wr_2053 ,           wr_2052 );
  nor g2627( wr_1029 , wr_1028 , wr_1000 );
  nor g2628( wr_1528 , wr_1527 , wr_718  );
  not g2629( G391    ,           wr_1552 );
  nor g2630( wr_744  , wr_743  , wr_617  );
  not g2631( wr_2796 ,           wr_2795 );
  not g2632( wr_2974 ,           wr_2973 );
  not g2633( wr_3117 ,           wr_3116 );
  not g2634( wr_3294 ,           wr_3293 );
  nor g2635( wr_2734 , wr_2733 , wr_2732 );
  nor g2636( wr_2799 , wr_2795 , wr_2798 );
  nor g2637( wr_2921 , wr_2920 , wr_2919 );
  nor g2638( wr_2977 , wr_2973 , wr_2976 );
  nor g2639( wr_3056 , wr_3055 , wr_3054 );
  nor g2640( wr_3120 , wr_3116 , wr_3119 );
  nor g2641( wr_3241 , wr_3240 , wr_3239 );
  nor g2642( wr_3297 , wr_3293 , wr_3296 );
  nor g2643( wr_1497 , wr_1469 , wr_743  );
  nor g2644( wr_363  , wr_362  , wr_288  );
  nor g2645( wr_567  , wr_566  , wr_489  );
  nor g2646( wr_2296 , wr_2295 , wr_667  );
  not g2647( wr_2836 ,           wr_2835 );
  not g2648( wr_3157 ,           wr_3156 );
  not g2649( wr_3334 ,           wr_3333 );
  not g2650( wr_1580 ,           wr_743  );
  nor g2651( wr_2838 , wr_2835 , wr_2541 );
  nor g2652( wr_3159 , wr_3156 , wr_2696 );
  nor g2653( wr_3336 , wr_3333 , wr_1622 );
  nor g2654( wr_2869 , wr_2868 , wr_2867 );
  nor g2655( wr_3190 , wr_3189 , wr_3188 );
  nor g2656( wr_3367 , wr_3366 , wr_3365 );
  nor g2657( wr_1440 , wr_1439 , wr_362  );
  nor g2658( wr_1459 , wr_1458 , wr_566  );
  nor g2659( wr_2334 , wr_2333 , wr_1479 );
  nor g2660( wr_1412 , wr_1411 , wr_1269 );
  nor g2661( wr_989  , wr_988  , wr_902  );
  nor g2662( wr_2262 , wr_2261 , wr_1334 );
  not g2663( wr_2327 ,           wr_403  );
  not g2664( wr_2499 ,           wr_362  );
  not g2665( wr_2654 ,           wr_566  );
  nor g2666( wr_687  , wr_686  , wr_164  );
  nor g2667( wr_1211 , wr_1210 , wr_1123 );
  nor g2668( wr_1355 , wr_1354 , wr_1335 );
  nor g2669( wr_1494 , wr_1493 , wr_164  );
  not g2670( wr_2313 ,           wr_1411 );
  nor g2671( wr_1842 , wr_1841 , wr_1688 );
  nor g2672( wr_2253 , wr_2252 , wr_2103 );
  nor g2673( wr_2054 , wr_2053 , wr_1892 );
  nor g2674( wr_404  , wr_403  , wr_183  );
  nor g2675( wr_1030 , wr_1029 , wr_767  );
  not g2676( wr_2255 ,           wr_1029 );
  not g2677( wr_2311 ,           wr_1210 );
  not g2678( wr_1529 ,           wr_1528 );
  nor g2679( wr_1532 , wr_1528 , wr_1531 );
  nor g2680( wr_745  , wr_744  , wr_711  );
  nor g2681( wr_2797 , wr_2796 , wr_2775 );
  nor g2682( wr_2975 , wr_2974 , wr_2953 );
  nor g2683( wr_3118 , wr_3117 , wr_3096 );
  nor g2684( wr_3295 , wr_3294 , wr_3273 );
  not g2685( wr_2735 ,           wr_2734 );
  not g2686( wr_2922 ,           wr_2921 );
  not g2687( wr_3057 ,           wr_3056 );
  not g2688( wr_3242 ,           wr_3241 );
  nor g2689( wr_1498 , wr_1497 , wr_711  );
  nor g2690( wr_2737 , wr_2734 , wr_2287 );
  nor g2691( wr_2924 , wr_2921 , wr_2307 );
  nor g2692( wr_3059 , wr_3056 , wr_2563 );
  nor g2693( wr_3244 , wr_3241 , wr_165  );
  nor g2694( wr_364  , wr_363  , wr_278  );
  nor g2695( wr_568  , wr_567  , wr_478  );
  nor g2696( wr_2837 , wr_2836 , wr_253  );
  nor g2697( wr_3158 , wr_3157 , wr_450  );
  nor g2698( wr_3335 , wr_3334 , wr_611  );
  nor g2699( wr_1582 , wr_1581 , wr_1580 );
  not g2700( wr_2870 ,           wr_2869 );
  not g2701( wr_3191 ,           wr_3190 );
  not g2702( wr_3368 ,           wr_3367 );
  nor g2703( wr_1441 , wr_1440 , wr_278  );
  nor g2704( wr_1460 , wr_1459 , wr_478  );
  nor g2705( wr_2872 , wr_2869 , wr_2494 );
  nor g2706( wr_3193 , wr_3190 , wr_2649 );
  nor g2707( wr_3370 , wr_3367 , wr_1575 );
  nor g2708( wr_1413 , wr_1412 , wr_1379 );
  nor g2709( wr_3080 , wr_3079 , wr_1580 );
  nor g2710( wr_990  , wr_989  , wr_892  );
  nor g2711( wr_2881 , wr_1449 , wr_2499 );
  nor g2712( wr_3017 , wr_1430 , wr_2327 );
  nor g2713( wr_3202 , wr_1486 , wr_2654 );
  nor g2714( wr_3379 , wr_1476 , wr_1580 );
  not g2715( wr_688  ,           wr_687  );
  nor g2716( wr_1212 , wr_1211 , wr_1112 );
  not g2717( wr_1356 ,           wr_1355 );
  not g2718( wr_1495 ,           wr_1494 );
  nor g2719( wr_2315 , wr_2314 , wr_2313 );
  not g2720( G412    ,           wr_1842 );
  not g2721( G416    ,           wr_2253 );
  not g2722( G414    ,           wr_2054 );
  nor g2723( wr_405  , wr_404  , wr_371  );
  nor g2724( wr_1031 , wr_1030 , wr_997  );
  nor g2725( wr_1530 , wr_1529 , wr_657  );
  nor g2726( wr_2297 , wr_745  , wr_421  );
  nor g2727( wr_2800 , wr_2799 , wr_2797 );
  nor g2728( wr_2978 , wr_2977 , wr_2975 );
  nor g2729( wr_3121 , wr_3120 , wr_3118 );
  nor g2730( wr_3298 , wr_3297 , wr_3295 );
  nor g2731( wr_2736 , wr_2735 , wr_411  );
  nor g2732( wr_2923 , wr_2922 , wr_194  );
  nor g2733( wr_3058 , wr_3057 , wr_672  );
  nor g2734( wr_3243 , wr_3242 , wr_162  );
  nor g2735( wr_2335 , wr_1498 , wr_1452 );
  not g2736( wr_2278 ,           wr_568  );
  not g2737( wr_2291 ,           wr_364  );
  nor g2738( wr_2839 , wr_2838 , wr_2837 );
  nor g2739( wr_3160 , wr_3159 , wr_3158 );
  nor g2740( wr_3337 , wr_3336 , wr_3335 );
  not g2741( wr_1583 ,           wr_1582 );
  nor g2742( wr_2277 , wr_745  , wr_682  );
  nor g2743( wr_2290 , wr_568  , wr_421  );
  nor g2744( wr_2559 , wr_2558 , wr_1582 );
  nor g2745( wr_2871 , wr_2870 , wr_239  );
  nor g2746( wr_3192 , wr_3191 , wr_431  );
  nor g2747( wr_3369 , wr_3368 , wr_601  );
  not g2748( wr_2329 ,           wr_1441 );
  not g2749( wr_2757 ,           wr_1460 );
  nor g2750( wr_2263 , wr_1413 , wr_1047 );
  not g2751( wr_3082 ,           wr_3080 );
  nor g2752( wr_2328 , wr_1460 , wr_1452 );
  nor g2753( wr_2756 , wr_1498 , wr_1489 );
  nor g2754( wr_3081 , wr_3080 , wr_3078 );
  nor g2755( wr_746  , wr_745  , wr_684  );
  nor g2756( wr_1414 , wr_1413 , wr_1352 );
  nor g2757( wr_1499 , wr_1498 , wr_1491 );
  not g2758( wr_2257 ,           wr_990  );
  not g2759( wr_2885 ,           wr_2881 );
  not g2760( wr_3021 ,           wr_3017 );
  not g2761( wr_3206 ,           wr_3202 );
  not g2762( wr_3383 ,           wr_3379 );
  nor g2763( wr_569  , wr_568  , wr_232  );
  nor g2764( wr_689  , wr_688  , wr_667  );
  nor g2765( wr_1213 , wr_1212 , wr_830  );
  nor g2766( wr_1357 , wr_1356 , wr_1334 );
  nor g2767( wr_1461 , wr_1460 , wr_1433 );
  nor g2768( wr_1496 , wr_1495 , wr_1479 );
  not g2769( wr_2317 ,           wr_2315 );
  nor g2770( wr_2256 , wr_1212 , wr_1047 );
  nor g2771( wr_2316 , wr_2315 , wr_2312 );
  nor g2772( wr_2475 , G416    , G412    );
  not g2773( wr_406  ,           wr_405  );
  not g2774( wr_1032 ,           wr_1031 );
  nor g2775( wr_365  , wr_364  , wr_232  );
  nor g2776( wr_991  , wr_990  , wr_830  );
  nor g2777( wr_1442 , wr_1441 , wr_1433 );
  nor g2778( wr_1600 , wr_1599 , wr_1582 );
  nor g2779( wr_1619 , wr_1618 , wr_1582 );
  nor g2780( wr_1632 , wr_1631 , wr_1582 );
  nor g2781( wr_1636 , wr_1582 , wr_1635 );
  nor g2782( wr_1533 , wr_1532 , wr_1530 );
  not g2783( wr_2298 ,           wr_2297 );
  not g2784( wr_2801 ,           wr_2800 );
  not g2785( wr_2979 ,           wr_2978 );
  not g2786( wr_3122 ,           wr_3121 );
  not g2787( wr_3299 ,           wr_3298 );
  nor g2788( wr_2738 , wr_2737 , wr_2736 );
  nor g2789( wr_2803 , wr_2800 , wr_2287 );
  nor g2790( wr_2925 , wr_2924 , wr_2923 );
  nor g2791( wr_2981 , wr_2978 , wr_2307 );
  nor g2792( wr_3060 , wr_3059 , wr_3058 );
  nor g2793( wr_3124 , wr_3121 , wr_2563 );
  nor g2794( wr_3245 , wr_3244 , wr_3243 );
  nor g2795( wr_3301 , wr_3298 , wr_165  );
  not g2796( wr_2336 ,           wr_2335 );
  nor g2797( wr_2282 , wr_2281 , wr_2278 );
  not g2798( wr_2840 ,           wr_2839 );
  not g2799( wr_3161 ,           wr_3160 );
  not g2800( wr_3338 ,           wr_3337 );
  nor g2801( wr_2557 , wr_1583 , wr_710  );
  nor g2802( wr_2842 , wr_2839 , wr_2494 );
  nor g2803( wr_3163 , wr_3160 , wr_2649 );
  nor g2804( wr_3340 , wr_3337 , wr_1575 );
  nor g2805( wr_2873 , wr_2872 , wr_2871 );
  nor g2806( wr_3194 , wr_3193 , wr_3192 );
  nor g2807( wr_3371 , wr_3370 , wr_3369 );
  nor g2808( wr_2761 , wr_2760 , wr_2757 );
  not g2809( wr_2264 ,           wr_2263 );
  nor g2810( wr_3083 , wr_3082 , wr_710  );
  not g2811( wr_747  ,           wr_746  );
  not g2812( wr_1415 ,           wr_1414 );
  not g2813( wr_1500 ,           wr_1499 );
  not g2814( wr_570  ,           wr_569  );
  not g2815( wr_1214 ,           wr_1213 );
  not g2816( wr_1462 ,           wr_1461 );
  nor g2817( wr_2318 , wr_2317 , wr_1378 );
  not g2818( wr_2476 ,           wr_2475 );
  nor g2819( wr_1584 , wr_1583 , wr_1579 );
  nor g2820( wr_1610 , wr_1609 , wr_1583 );
  nor g2821( wr_1625 , wr_1624 , wr_1583 );
  nor g2822( wr_1634 , wr_1583 , wr_581  );
  not g2823( G388    ,           wr_1533 );
  nor g2824( wr_2299 , wr_2298 , wr_682  );
  nor g2825( wr_2802 , wr_2801 , wr_411  );
  nor g2826( wr_2980 , wr_2979 , wr_194  );
  nor g2827( wr_3123 , wr_3122 , wr_672  );
  nor g2828( wr_3300 , wr_3299 , wr_162  );
  not g2829( wr_2739 ,           wr_2738 );
  not g2830( wr_2926 ,           wr_2925 );
  not g2831( wr_3061 ,           wr_3060 );
  not g2832( wr_3246 ,           wr_3245 );
  nor g2833( wr_2337 , wr_2336 , wr_1489 );
  nor g2834( wr_2741 , wr_2738 , wr_2408 );
  nor g2835( wr_2928 , wr_2925 , wr_2470 );
  nor g2836( wr_3063 , wr_3060 , wr_2642 );
  nor g2837( wr_3248 , wr_3245 , wr_1568 );
  not g2838( wr_2283 ,           wr_2282 );
  nor g2839( wr_2841 , wr_2840 , wr_239  );
  nor g2840( wr_3162 , wr_3161 , wr_431  );
  nor g2841( wr_3339 , wr_3338 , wr_601  );
  nor g2842( wr_2560 , wr_2559 , wr_2557 );
  not g2843( wr_2874 ,           wr_2873 );
  not g2844( wr_3195 ,           wr_3194 );
  not g2845( wr_3372 ,           wr_3371 );
  not g2846( wr_2762 ,           wr_2761 );
  nor g2847( wr_2876 , wr_2873 , wr_2524 );
  nor g2848( wr_3197 , wr_3194 , wr_2679 );
  nor g2849( wr_3374 , wr_3371 , wr_1605 );
  nor g2850( wr_2265 , wr_2264 , wr_1350 );
  nor g2851( wr_3084 , wr_3083 , wr_3081 );
  nor g2852( wr_748  , wr_747  , wr_682  );
  nor g2853( wr_1416 , wr_1415 , wr_1350 );
  nor g2854( wr_1501 , wr_1500 , wr_1489 );
  nor g2855( wr_571  , wr_570  , wr_421  );
  nor g2856( wr_1215 , wr_1214 , wr_1047 );
  nor g2857( wr_1463 , wr_1462 , wr_1452 );
  nor g2858( wr_2319 , wr_2318 , wr_2316 );
  nor g2859( wr_2477 , wr_2476 , G414    );
  nor g2860( wr_1601 , wr_1600 , wr_1584 );
  nor g2861( wr_1620 , wr_1619 , wr_1610 );
  nor g2862( wr_1633 , wr_1632 , wr_1625 );
  nor g2863( wr_1637 , wr_1636 , wr_1634 );
  nor g2864( wr_2300 , wr_2299 , wr_2296 );
  nor g2865( wr_2804 , wr_2803 , wr_2802 );
  nor g2866( wr_2982 , wr_2981 , wr_2980 );
  nor g2867( wr_3125 , wr_3124 , wr_3123 );
  nor g2868( wr_3302 , wr_3301 , wr_3300 );
  nor g2869( wr_2740 , wr_2739 , wr_334  );
  nor g2870( wr_2927 , wr_2926 , wr_215  );
  nor g2871( wr_3062 , wr_3061 , wr_538  );
  nor g2872( wr_3247 , wr_3246 , wr_647  );
  nor g2873( wr_2338 , wr_2337 , wr_2334 );
  nor g2874( wr_2284 , wr_2283 , wr_2277 );
  nor g2875( wr_2843 , wr_2842 , wr_2841 );
  nor g2876( wr_3164 , wr_3163 , wr_3162 );
  nor g2877( wr_3341 , wr_3340 , wr_3339 );
  nor g2878( wr_2590 , wr_2589 , wr_2560 );
  nor g2879( wr_2875 , wr_2874 , wr_257  );
  nor g2880( wr_3196 , wr_3195 , wr_455  );
  nor g2881( wr_3373 , wr_3372 , wr_591  );
  nor g2882( wr_2611 , wr_2610 , wr_2560 );
  nor g2883( wr_2763 , wr_2762 , wr_2756 );
  nor g2884( wr_2266 , wr_2265 , wr_2262 );
  nor g2885( wr_2627 , wr_2560 , wr_538  );
  not g2886( wr_3085 ,           wr_3084 );
  nor g2887( wr_749  , wr_748  , wr_689  );
  nor g2888( wr_1417 , wr_1416 , wr_1357 );
  nor g2889( wr_1502 , wr_1501 , wr_1496 );
  nor g2890( wr_2320 , wr_2319 , wr_1348 );
  nor g2891( wr_2638 , wr_2560 , wr_672  );
  nor g2892( wr_2655 , wr_2560 , wr_680  );
  not g2893( wr_2478 ,           wr_2477 );
  not g2894( wr_2561 ,           wr_2560 );
  nor g2895( wr_2564 , wr_2560 , wr_2563 );
  not g2896( G376    ,           wr_1601 );
  not g2897( G379    ,           wr_1620 );
  not g2898( G382    ,           wr_1633 );
  not g2899( G385    ,           wr_1637 );
  not g2900( wr_2301 ,           wr_2300 );
  not g2901( wr_2805 ,           wr_2804 );
  not g2902( wr_2983 ,           wr_2982 );
  not g2903( wr_3126 ,           wr_3125 );
  not g2904( wr_3303 ,           wr_3302 );
  nor g2905( wr_2742 , wr_2741 , wr_2740 );
  nor g2906( wr_2807 , wr_2804 , wr_2408 );
  nor g2907( wr_2929 , wr_2928 , wr_2927 );
  nor g2908( wr_2985 , wr_2982 , wr_2470 );
  nor g2909( wr_3064 , wr_3063 , wr_3062 );
  nor g2910( wr_3128 , wr_3125 , wr_2642 );
  nor g2911( wr_3249 , wr_3248 , wr_3247 );
  nor g2912( wr_3305 , wr_3302 , wr_1568 );
  not g2913( wr_2339 ,           wr_2338 );
  nor g2914( wr_2356 , wr_2355 , wr_2284 );
  not g2915( wr_2844 ,           wr_2843 );
  not g2916( wr_3165 ,           wr_3164 );
  not g2917( wr_3342 ,           wr_3341 );
  not g2918( wr_2591 ,           wr_2590 );
  nor g2919( wr_2846 , wr_2843 , wr_2524 );
  nor g2920( wr_3167 , wr_3164 , wr_2679 );
  nor g2921( wr_3344 , wr_3341 , wr_1605 );
  nor g2922( wr_2377 , wr_2376 , wr_2284 );
  nor g2923( wr_2877 , wr_2876 , wr_2875 );
  nor g2924( wr_3198 , wr_3197 , wr_3196 );
  nor g2925( wr_3375 , wr_3374 , wr_3373 );
  not g2926( wr_2612 ,           wr_2611 );
  not g2927( wr_2267 ,           wr_2266 );
  nor g2928( wr_2393 , wr_2284 , wr_334  );
  not g2929( wr_2764 ,           wr_2763 );
  not g2930( wr_2628 ,           wr_2627 );
  not g2931( wr_750  ,           wr_749  );
  not g2932( wr_1418 ,           wr_1417 );
  not g2933( wr_1503 ,           wr_1502 );
  nor g2934( wr_2404 , wr_2284 , wr_411  );
  nor g2935( wr_2500 , wr_2284 , wr_419  );
  nor g2936( wr_2321 , wr_2320 , wr_2311 );
  nor g2937( wr_2639 , wr_2638 , wr_544  );
  nor g2938( wr_2656 , wr_2655 , wr_2654 );
  not g2939( wr_2285 ,           wr_2284 );
  nor g2940( wr_2481 , wr_2480 , wr_2478 );
  nor g2941( wr_2288 , wr_2284 , wr_2287 );
  nor g2942( wr_2562 , wr_2561 , wr_672  );
  nor g2943( wr_2302 , wr_2301 , wr_2291 );
  nor g2944( wr_2806 , wr_2805 , wr_334  );
  nor g2945( wr_2984 , wr_2983 , wr_215  );
  nor g2946( wr_3127 , wr_3126 , wr_538  );
  nor g2947( wr_3304 , wr_3303 , wr_647  );
  not g2948( wr_2743 ,           wr_2742 );
  not g2949( wr_2930 ,           wr_2929 );
  not g2950( wr_3065 ,           wr_3064 );
  not g2951( wr_3250 ,           wr_3249 );
  nor g2952( wr_2340 , wr_2339 , wr_2329 );
  nor g2953( wr_2745 , wr_2742 , wr_2371 );
  nor g2954( wr_2932 , wr_2929 , wr_2433 );
  nor g2955( wr_3067 , wr_3064 , wr_2605 );
  nor g2956( wr_3252 , wr_3249 , wr_1531 );
  not g2957( wr_2357 ,           wr_2356 );
  nor g2958( wr_2845 , wr_2844 , wr_257  );
  nor g2959( wr_3166 , wr_3165 , wr_455  );
  nor g2960( wr_3343 , wr_3342 , wr_591  );
  nor g2961( wr_2592 , wr_2591 , wr_672  );
  not g2962( wr_2378 ,           wr_2377 );
  nor g2963( wr_2886 , wr_2877 , wr_2763 );
  nor g2964( wr_3207 , wr_3198 , wr_3084 );
  nor g2965( wr_3384 , wr_3375 , wr_164  );
  nor g2966( wr_2613 , wr_2612 , wr_672  );
  nor g2967( wr_2268 , wr_2267 , wr_2257 );
  not g2968( wr_2394 ,           wr_2393 );
  nor g2969( wr_2878 , wr_2877 , wr_2764 );
  nor g2970( wr_3199 , wr_3198 , wr_3085 );
  nor g2971( wr_3376 , wr_3375 , G4526   );
  nor g2972( wr_2629 , wr_2628 , wr_672  );
  nor g2973( wr_751  , wr_750  , wr_571  );
  nor g2974( wr_1419 , wr_1418 , wr_1215 );
  nor g2975( wr_1504 , wr_1503 , wr_1463 );
  nor g2976( wr_2405 , wr_2404 , wr_340  );
  nor g2977( wr_2501 , wr_2500 , wr_2499 );
  not g2978( wr_2323 ,           wr_2321 );
  not g2979( wr_2640 ,           wr_2639 );
  not g2980( wr_2657 ,           wr_2656 );
  nor g2981( wr_2286 , wr_2285 , wr_411  );
  nor g2982( wr_2322 , wr_2321 , wr_2310 );
  not g2983( wr_2482 ,           wr_2481 );
  nor g2984( wr_2643 , wr_2639 , wr_2642 );
  nor g2985( wr_2674 , wr_2673 , wr_2656 );
  nor g2986( wr_2693 , wr_2692 , wr_2656 );
  nor g2987( wr_2706 , wr_2705 , wr_2656 );
  nor g2988( wr_2710 , wr_2656 , wr_2709 );
  nor g2989( wr_2565 , wr_2564 , wr_2562 );
  not g2990( wr_2303 ,           wr_2302 );
  nor g2991( wr_2808 , wr_2807 , wr_2806 );
  nor g2992( wr_2986 , wr_2985 , wr_2984 );
  nor g2993( wr_3129 , wr_3128 , wr_3127 );
  nor g2994( wr_3306 , wr_3305 , wr_3304 );
  nor g2995( wr_2744 , wr_2743 , wr_295  );
  nor g2996( wr_2931 , wr_2930 , wr_222  );
  nor g2997( wr_3066 , wr_3065 , wr_499  );
  nor g2998( wr_3251 , wr_3250 , wr_657  );
  not g2999( wr_2341 ,           wr_2340 );
  nor g3000( wr_2358 , wr_2357 , wr_411  );
  nor g3001( wr_2847 , wr_2846 , wr_2845 );
  nor g3002( wr_3168 , wr_3167 , wr_3166 );
  nor g3003( wr_3345 , wr_3344 , wr_3343 );
  nor g3004( wr_2596 , wr_2595 , wr_2592 );
  nor g3005( wr_2379 , wr_2378 , wr_411  );
  not g3006( wr_2887 ,           wr_2886 );
  not g3007( wr_3208 ,           wr_3207 );
  not g3008( wr_3385 ,           wr_3384 );
  nor g3009( wr_2617 , wr_2616 , wr_2613 );
  not g3010( wr_2269 ,           wr_2268 );
  nor g3011( wr_2395 , wr_2394 , wr_411  );
  not g3012( wr_2879 ,           wr_2878 );
  not g3013( wr_3200 ,           wr_3199 );
  not g3014( wr_3377 ,           wr_3376 );
  nor g3015( wr_2630 , wr_2629 , wr_553  );
  not g3016( wr_752  ,           wr_751  );
  not g3017( wr_1420 ,           wr_1419 );
  not g3018( wr_1505 ,           wr_1504 );
  not g3019( wr_2406 ,           wr_2405 );
  not g3020( wr_2502 ,           wr_2501 );
  nor g3021( wr_2324 , wr_2323 , wr_1111 );
  nor g3022( wr_2409 , wr_2405 , wr_2408 );
  nor g3023( wr_2519 , wr_2518 , wr_2501 );
  nor g3024( wr_2538 , wr_2537 , wr_2501 );
  nor g3025( wr_2551 , wr_2550 , wr_2501 );
  nor g3026( wr_2555 , wr_2501 , wr_2554 );
  nor g3027( wr_2641 , wr_2640 , wr_538  );
  nor g3028( wr_2658 , wr_2657 , wr_2653 );
  nor g3029( wr_2684 , wr_2683 , wr_2657 );
  nor g3030( wr_2699 , wr_2698 , wr_2657 );
  nor g3031( wr_2708 , wr_2657 , wr_483  );
  nor g3032( wr_2289 , wr_2288 , wr_2286 );
  nor g3033( wr_2483 , wr_2482 , wr_2474 );
  not g3034( G344    ,           wr_2565 );
  nor g3035( wr_2304 , wr_2303 , wr_2290 );
  not g3036( wr_2809 ,           wr_2808 );
  not g3037( wr_2987 ,           wr_2986 );
  not g3038( wr_3130 ,           wr_3129 );
  not g3039( wr_3307 ,           wr_3306 );
  nor g3040( wr_2746 , wr_2745 , wr_2744 );
  nor g3041( wr_2811 , wr_2808 , wr_2371 );
  nor g3042( wr_2933 , wr_2932 , wr_2931 );
  nor g3043( wr_2989 , wr_2986 , wr_2433 );
  nor g3044( wr_3068 , wr_3067 , wr_3066 );
  nor g3045( wr_3132 , wr_3129 , wr_2605 );
  nor g3046( wr_3253 , wr_3252 , wr_3251 );
  nor g3047( wr_3309 , wr_3306 , wr_1531 );
  nor g3048( wr_2342 , wr_2341 , wr_2328 );
  nor g3049( wr_2362 , wr_2361 , wr_2358 );
  nor g3050( wr_2882 , wr_2847 , wr_2763 );
  nor g3051( wr_3203 , wr_3168 , wr_3084 );
  nor g3052( wr_3380 , wr_3345 , wr_164  );
  not g3053( wr_2597 ,           wr_2596 );
  nor g3054( wr_2383 , wr_2382 , wr_2379 );
  nor g3055( wr_2888 , wr_2887 , wr_2885 );
  nor g3056( wr_3209 , wr_3208 , wr_3206 );
  nor g3057( wr_3386 , wr_3385 , wr_3383 );
  not g3058( wr_2618 ,           wr_2617 );
  nor g3059( wr_2270 , wr_2269 , wr_2256 );
  nor g3060( wr_2396 , wr_2395 , wr_349  );
  nor g3061( wr_2848 , wr_2847 , wr_2764 );
  nor g3062( wr_2880 , wr_2879 , wr_2499 );
  nor g3063( wr_3169 , wr_3168 , wr_3085 );
  nor g3064( wr_3201 , wr_3200 , wr_2654 );
  nor g3065( wr_3346 , wr_3345 , G4526   );
  nor g3066( wr_3378 , wr_3377 , wr_1580 );
  not g3067( wr_2631 ,           wr_2630 );
  nor g3068( wr_753  , wr_752  , wr_406  );
  nor g3069( wr_1421 , wr_1420 , wr_1032 );
  nor g3070( wr_1506 , wr_1505 , wr_406  );
  nor g3071( wr_2407 , wr_2406 , wr_334  );
  nor g3072( wr_2503 , wr_2502 , wr_2498 );
  nor g3073( wr_2529 , wr_2528 , wr_2502 );
  nor g3074( wr_2544 , wr_2543 , wr_2502 );
  nor g3075( wr_2553 , wr_2502 , wr_282  );
  nor g3076( wr_2325 , wr_2324 , wr_2322 );
  nor g3077( wr_2644 , wr_2643 , wr_2641 );
  nor g3078( wr_2675 , wr_2674 , wr_2658 );
  nor g3079( wr_2694 , wr_2693 , wr_2684 );
  nor g3080( wr_2707 , wr_2706 , wr_2699 );
  nor g3081( wr_2711 , wr_2710 , wr_2708 );
  not g3082( G295    ,           wr_2289 );
  not g3083( G418    ,           wr_2483 );
  nor g3084( wr_2418 , wr_2417 , wr_2304 );
  nor g3085( wr_2810 , wr_2809 , wr_295  );
  nor g3086( wr_2988 , wr_2987 , wr_222  );
  nor g3087( wr_3131 , wr_3130 , wr_499  );
  nor g3088( wr_3308 , wr_3307 , wr_657  );
  nor g3089( wr_2439 , wr_2438 , wr_2304 );
  not g3090( wr_2747 ,           wr_2746 );
  not g3091( wr_2934 ,           wr_2933 );
  not g3092( wr_3069 ,           wr_3068 );
  not g3093( wr_3254 ,           wr_3253 );
  nor g3094( wr_2749 , wr_2746 , wr_2401 );
  nor g3095( wr_2936 , wr_2933 , wr_2463 );
  nor g3096( wr_3018 , wr_3005 , wr_2342 );
  nor g3097( wr_3022 , wr_3013 , wr_2342 );
  nor g3098( wr_3071 , wr_3068 , wr_2635 );
  nor g3099( wr_3256 , wr_3253 , wr_1561 );
  not g3100( wr_2363 ,           wr_2362 );
  nor g3101( wr_2455 , wr_2304 , wr_215  );
  not g3102( wr_2883 ,           wr_2882 );
  not g3103( wr_2898 ,           wr_2342 );
  not g3104( wr_3204 ,           wr_3203 );
  not g3105( wr_3381 ,           wr_3380 );
  nor g3106( wr_2598 , wr_2597 , wr_2585 );
  not g3107( wr_2384 ,           wr_2383 );
  nor g3108( wr_2619 , wr_2618 , wr_519  );
  nor g3109( wr_2271 , wr_2270 , wr_828  );
  nor g3110( wr_2343 , wr_2342 , wr_1431 );
  not g3111( wr_2397 ,           wr_2396 );
  nor g3112( wr_2466 , wr_2304 , wr_194  );
  nor g3113( wr_2484 , wr_2304 , wr_230  );
  not g3114( wr_2849 ,           wr_2848 );
  not g3115( wr_3170 ,           wr_3169 );
  not g3116( wr_3347 ,           wr_3346 );
  nor g3117( wr_2632 , wr_2631 , wr_2614 );
  not g3118( wr_2305 ,           wr_2304 );
  not g3119( wr_754  ,           wr_753  );
  not g3120( wr_1422 ,           wr_1421 );
  not g3121( wr_1507 ,           wr_1506 );
  nor g3122( wr_2308 , wr_2304 , wr_2307 );
  nor g3123( wr_2410 , wr_2409 , wr_2407 );
  nor g3124( wr_2520 , wr_2519 , wr_2503 );
  nor g3125( wr_2539 , wr_2538 , wr_2529 );
  nor g3126( wr_2552 , wr_2551 , wr_2544 );
  nor g3127( wr_2556 , wr_2555 , wr_2553 );
  not g3128( G252    ,           wr_2325 );
  not g3129( G368    ,           wr_2644 );
  not g3130( G347    ,           wr_2675 );
  not g3131( G350    ,           wr_2694 );
  not g3132( G353    ,           wr_2707 );
  not g3133( G356    ,           wr_2711 );
  not g3134( wr_2419 ,           wr_2418 );
  nor g3135( wr_2812 , wr_2811 , wr_2810 );
  nor g3136( wr_2990 , wr_2989 , wr_2988 );
  nor g3137( wr_3133 , wr_3132 , wr_3131 );
  nor g3138( wr_3310 , wr_3309 , wr_3308 );
  not g3139( wr_2440 ,           wr_2439 );
  nor g3140( wr_2748 , wr_2747 , wr_324  );
  nor g3141( wr_2935 , wr_2934 , wr_208  );
  nor g3142( wr_3070 , wr_3069 , wr_528  );
  nor g3143( wr_3255 , wr_3254 , wr_637  );
  not g3144( wr_3019 ,           wr_3018 );
  not g3145( wr_3023 ,           wr_3022 );
  nor g3146( wr_2364 , wr_2363 , wr_2351 );
  not g3147( wr_2456 ,           wr_2455 );
  nor g3148( wr_2884 , wr_2883 , wr_2881 );
  nor g3149( wr_3014 , wr_3013 , wr_2898 );
  nor g3150( wr_3205 , wr_3204 , wr_3202 );
  nor g3151( wr_3382 , wr_3381 , wr_3379 );
  not g3152( wr_2599 ,           wr_2598 );
  nor g3153( wr_2385 , wr_2384 , wr_315  );
  nor g3154( wr_3006 , wr_3005 , wr_2898 );
  not g3155( wr_2620 ,           wr_2619 );
  nor g3156( wr_2272 , wr_2271 , wr_2255 );
  nor g3157( wr_2344 , wr_2343 , wr_2327 );
  nor g3158( wr_2398 , wr_2397 , wr_2380 );
  nor g3159( wr_2467 , wr_2466 , wr_381  );
  nor g3160( wr_2485 , wr_2484 , wr_2327 );
  nor g3161( wr_2850 , wr_2849 , wr_362  );
  nor g3162( wr_3171 , wr_3170 , wr_566  );
  nor g3163( wr_3348 , wr_3347 , wr_743  );
  not g3164( wr_2633 ,           wr_2632 );
  nor g3165( wr_2306 , wr_2305 , wr_194  );
  nor g3166( wr_2636 , wr_2632 , wr_2635 );
  nor g3167( wr_755  , wr_754  , wr_365  );
  nor g3168( wr_1423 , wr_1422 , wr_991  );
  nor g3169( wr_1508 , wr_1507 , wr_1442 );
  not g3170( G319    ,           wr_2410 );
  not g3171( G298    ,           wr_2520 );
  not g3172( G301    ,           wr_2539 );
  not g3173( G304    ,           wr_2552 );
  not g3174( G307    ,           wr_2556 );
  nor g3175( wr_2420 , wr_2419 , wr_194  );
  not g3176( wr_2813 ,           wr_2812 );
  not g3177( wr_2991 ,           wr_2990 );
  not g3178( wr_3134 ,           wr_3133 );
  not g3179( wr_3311 ,           wr_3310 );
  nor g3180( wr_2441 , wr_2440 , wr_194  );
  nor g3181( wr_2750 , wr_2749 , wr_2748 );
  nor g3182( wr_2815 , wr_2812 , wr_2401 );
  nor g3183( wr_2937 , wr_2936 , wr_2935 );
  nor g3184( wr_2993 , wr_2990 , wr_2463 );
  nor g3185( wr_3072 , wr_3071 , wr_3070 );
  nor g3186( wr_3136 , wr_3133 , wr_2635 );
  nor g3187( wr_3257 , wr_3256 , wr_3255 );
  nor g3188( wr_3313 , wr_3310 , wr_1561 );
  nor g3189( wr_3020 , wr_3019 , wr_3017 );
  nor g3190( wr_3024 , wr_3023 , wr_3021 );
  not g3191( wr_2365 ,           wr_2364 );
  nor g3192( wr_2457 , wr_2456 , wr_194  );
  nor g3193( wr_2889 , wr_2888 , wr_2884 );
  not g3194( wr_3015 ,           wr_3014 );
  nor g3195( wr_3210 , wr_3209 , wr_3205 );
  nor g3196( wr_3387 , wr_3386 , wr_3382 );
  nor g3197( wr_2600 , wr_2599 , wr_505  );
  not g3198( wr_2386 ,           wr_2385 );
  not g3199( wr_3007 ,           wr_3006 );
  nor g3200( wr_2621 , wr_2620 , wr_2608 );
  not g3201( wr_2274 ,           wr_2272 );
  not g3202( wr_2346 ,           wr_2344 );
  not g3203( wr_2399 ,           wr_2398 );
  not g3204( wr_2468 ,           wr_2467 );
  not g3205( wr_2486 ,           wr_2485 );
  nor g3206( wr_2273 , wr_2272 , wr_2254 );
  nor g3207( wr_2345 , wr_2344 , wr_2326 );
  nor g3208( wr_2402 , wr_2398 , wr_2401 );
  nor g3209( wr_2471 , wr_2467 , wr_2470 );
  nor g3210( wr_2488 , wr_2485 , wr_2326 );
  nor g3211( wr_2577 , wr_2576 , wr_2485 );
  nor g3212( wr_2581 , wr_2485 , wr_2580 );
  nor g3213( wr_2634 , wr_2633 , wr_528  );
  nor g3214( wr_2309 , wr_2308 , wr_2306 );
  not g3215( G246    ,           wr_755  );
  not g3216( G258    ,           wr_1423 );
  not g3217( G270    ,           wr_1508 );
  not g3218( G264    ,           wr_1423 );
  nor g3219( wr_2424 , wr_2423 , wr_2420 );
  nor g3220( wr_2814 , wr_2813 , wr_324  );
  nor g3221( wr_2992 , wr_2991 , wr_208  );
  nor g3222( wr_3135 , wr_3134 , wr_528  );
  nor g3223( wr_3312 , wr_3311 , wr_637  );
  nor g3224( wr_2445 , wr_2444 , wr_2441 );
  not g3225( wr_2751 ,           wr_2750 );
  not g3226( wr_2938 ,           wr_2937 );
  not g3227( wr_3073 ,           wr_3072 );
  not g3228( wr_3258 ,           wr_3257 );
  nor g3229( wr_2753 , wr_2750 , wr_2390 );
  nor g3230( wr_2940 , wr_2937 , wr_2452 );
  nor g3231( wr_3025 , wr_3024 , wr_3020 );
  nor g3232( wr_3075 , wr_3072 , wr_2624 );
  nor g3233( wr_3260 , wr_3257 , wr_1550 );
  nor g3234( wr_2366 , wr_2365 , wr_301  );
  nor g3235( wr_2458 , wr_2457 , wr_390  );
  not g3236( wr_2890 ,           wr_2889 );
  nor g3237( wr_3016 , wr_3015 , wr_2327 );
  not g3238( wr_3211 ,           wr_3210 );
  not g3239( wr_3388 ,           wr_3387 );
  not g3240( wr_2601 ,           wr_2600 );
  nor g3241( wr_2387 , wr_2386 , wr_2374 );
  nor g3242( wr_3008 , wr_3007 , wr_403  );
  not g3243( wr_2622 ,           wr_2621 );
  nor g3244( wr_2275 , wr_2274 , wr_996  );
  nor g3245( wr_2347 , wr_2346 , wr_370  );
  nor g3246( wr_2400 , wr_2399 , wr_324  );
  nor g3247( wr_2469 , wr_2468 , wr_215  );
  nor g3248( wr_2487 , wr_2486 , wr_370  );
  nor g3249( wr_2570 , wr_2569 , wr_2486 );
  nor g3250( wr_2579 , wr_2486 , wr_175  );
  nor g3251( wr_2625 , wr_2621 , wr_2624 );
  nor g3252( wr_2637 , wr_2636 , wr_2634 );
  not g3253( G324    ,           wr_2309 );
  not g3254( wr_2425 ,           wr_2424 );
  nor g3255( wr_2816 , wr_2815 , wr_2814 );
  nor g3256( wr_2994 , wr_2993 , wr_2992 );
  nor g3257( wr_3137 , wr_3136 , wr_3135 );
  nor g3258( wr_3314 , wr_3313 , wr_3312 );
  not g3259( wr_2446 ,           wr_2445 );
  nor g3260( wr_2752 , wr_2751 , wr_309  );
  nor g3261( wr_2939 , wr_2938 , wr_201  );
  nor g3262( wr_3074 , wr_3073 , wr_513  );
  nor g3263( wr_3259 , wr_3258 , wr_627  );
  not g3264( wr_3026 ,           wr_3025 );
  not g3265( wr_2367 ,           wr_2366 );
  not g3266( wr_2459 ,           wr_2458 );
  nor g3267( wr_2891 , wr_2890 , wr_2880 );
  nor g3268( wr_3212 , wr_3211 , wr_3201 );
  nor g3269( wr_3389 , wr_3388 , wr_3378 );
  nor g3270( wr_2602 , wr_2601 , wr_521  );
  not g3271( wr_2388 ,           wr_2387 );
  nor g3272( wr_2391 , wr_2387 , wr_2390 );
  nor g3273( wr_2623 , wr_2622 , wr_513  );
  nor g3274( wr_2276 , wr_2275 , wr_2273 );
  nor g3275( wr_2348 , wr_2347 , wr_2345 );
  nor g3276( wr_2403 , wr_2402 , wr_2400 );
  nor g3277( wr_2472 , wr_2471 , wr_2469 );
  nor g3278( wr_2489 , wr_2488 , wr_2487 );
  nor g3279( wr_2578 , wr_2577 , wr_2570 );
  nor g3280( wr_2582 , wr_2581 , wr_2579 );
  not g3281( G365    ,           wr_2637 );
  nor g3282( wr_2426 , wr_2425 , wr_2413 );
  not g3283( wr_2817 ,           wr_2816 );
  not g3284( wr_2995 ,           wr_2994 );
  not g3285( wr_3138 ,           wr_3137 );
  not g3286( wr_3315 ,           wr_3314 );
  nor g3287( wr_2447 , wr_2446 , wr_376  );
  nor g3288( wr_2754 , wr_2753 , wr_2752 );
  nor g3289( wr_2819 , wr_2816 , wr_2390 );
  nor g3290( wr_2941 , wr_2940 , wr_2939 );
  nor g3291( wr_2997 , wr_2994 , wr_2452 );
  nor g3292( wr_3076 , wr_3075 , wr_3074 );
  nor g3293( wr_3140 , wr_3137 , wr_2624 );
  nor g3294( wr_3261 , wr_3260 , wr_3259 );
  nor g3295( wr_3317 , wr_3314 , wr_1550 );
  nor g3296( wr_3027 , wr_3026 , wr_3016 );
  nor g3297( wr_2368 , wr_2367 , wr_317  );
  nor g3298( wr_2460 , wr_2459 , wr_2442 );
  not g3299( wr_2892 ,           wr_2891 );
  not g3300( wr_3213 ,           wr_3212 );
  not g3301( wr_3390 ,           wr_3389 );
  not g3302( wr_2603 ,           wr_2602 );
  nor g3303( wr_2389 , wr_2388 , wr_309  );
  nor g3304( wr_2606 , wr_2602 , wr_2605 );
  nor g3305( wr_2626 , wr_2625 , wr_2623 );
  not g3306( G249    ,           wr_2276 );
  not g3307( G276    ,           wr_2348 );
  not g3308( G316    ,           wr_2403 );
  not g3309( G336    ,           wr_2472 );
  not g3310( G273    ,           wr_2489 );
  not g3311( G422    ,           wr_2578 );
  not g3312( G419    ,           wr_2582 );
  not g3313( G469    ,           wr_2578 );
  not g3314( G471    ,           wr_2582 );
  not g3315( wr_2427 ,           wr_2426 );
  nor g3316( wr_2818 , wr_2817 , wr_309  );
  nor g3317( wr_2996 , wr_2995 , wr_201  );
  nor g3318( wr_3139 , wr_3138 , wr_513  );
  nor g3319( wr_3316 , wr_3315 , wr_627  );
  not g3320( wr_2448 ,           wr_2447 );
  not g3321( wr_2755 ,           wr_2754 );
  not g3322( wr_2942 ,           wr_2941 );
  not g3323( wr_3077 ,           wr_3076 );
  not g3324( wr_3262 ,           wr_3261 );
  not g3325( wr_3028 ,           wr_3027 );
  not g3326( wr_2369 ,           wr_2368 );
  not g3327( wr_2461 ,           wr_2460 );
  nor g3328( wr_2893 , wr_2892 , wr_2850 );
  nor g3329( wr_3214 , wr_3213 , wr_3171 );
  nor g3330( wr_3391 , wr_3390 , wr_3348 );
  nor g3331( wr_2372 , wr_2368 , wr_2371 );
  nor g3332( wr_2464 , wr_2460 , wr_2463 );
  nor g3333( wr_2604 , wr_2603 , wr_499  );
  nor g3334( wr_2392 , wr_2391 , wr_2389 );
  not g3335( G362    ,           wr_2626 );
  nor g3336( wr_2428 , wr_2427 , wr_372  );
  nor g3337( wr_2820 , wr_2819 , wr_2818 );
  nor g3338( wr_2998 , wr_2997 , wr_2996 );
  nor g3339( wr_3141 , wr_3140 , wr_3139 );
  nor g3340( wr_3318 , wr_3317 , wr_3316 );
  nor g3341( wr_2449 , wr_2448 , wr_2436 );
  nor g3342( wr_2765 , wr_2764 , wr_2755 );
  nor g3343( wr_2943 , wr_2942 , wr_2898 );
  nor g3344( wr_3086 , wr_3085 , wr_3077 );
  nor g3345( wr_3263 , wr_3262 , G4526   );
  nor g3346( wr_3029 , wr_3028 , wr_3008 );
  nor g3347( wr_2370 , wr_2369 , wr_295  );
  nor g3348( wr_2462 , wr_2461 , wr_208  );
  not g3349( wr_2894 ,           wr_2893 );
  not g3350( wr_3215 ,           wr_3214 );
  not g3351( wr_3392 ,           wr_3391 );
  nor g3352( wr_2607 , wr_2606 , wr_2604 );
  not g3353( G313    ,           wr_2392 );
  not g3354( wr_2429 ,           wr_2428 );
  nor g3355( wr_2821 , wr_2820 , wr_2763 );
  nor g3356( wr_2999 , wr_2998 , wr_2342 );
  nor g3357( wr_3142 , wr_3141 , wr_3084 );
  nor g3358( wr_3319 , wr_3318 , wr_164  );
  not g3359( wr_2450 ,           wr_2449 );
  nor g3360( wr_2453 , wr_2449 , wr_2452 );
  not g3361( wr_3030 ,           wr_3029 );
  nor g3362( wr_2373 , wr_2372 , wr_2370 );
  nor g3363( wr_2465 , wr_2464 , wr_2462 );
  not g3364( G359    ,           wr_2607 );
  nor g3365( wr_2430 , wr_2429 , wr_378  );
  nor g3366( wr_2822 , wr_2821 , wr_2765 );
  nor g3367( wr_3000 , wr_2999 , wr_2943 );
  nor g3368( wr_3143 , wr_3142 , wr_3086 );
  nor g3369( wr_3320 , wr_3319 , wr_3263 );
  nor g3370( wr_2451 , wr_2450 , wr_201  );
  not g3371( G310    ,           wr_2373 );
  not g3372( G333    ,           wr_2465 );
  not g3373( wr_2431 ,           wr_2430 );
  nor g3374( wr_2434 , wr_2430 , wr_2433 );
  not g3375( wr_2896 ,           wr_2822 );
  not g3376( wr_3032 ,           wr_3000 );
  not g3377( wr_3217 ,           wr_3143 );
  not g3378( wr_3394 ,           wr_3320 );
  nor g3379( wr_2454 , wr_2453 , wr_2451 );
  nor g3380( wr_2895 , wr_2894 , wr_2822 );
  nor g3381( wr_3031 , wr_3030 , wr_3000 );
  nor g3382( wr_3216 , wr_3215 , wr_3143 );
  nor g3383( wr_3393 , wr_3392 , wr_3320 );
  nor g3384( wr_2432 , wr_2431 , wr_222  );
  nor g3385( wr_2897 , wr_2893 , wr_2896 );
  nor g3386( wr_3033 , wr_3029 , wr_3032 );
  nor g3387( wr_3218 , wr_3214 , wr_3217 );
  nor g3388( wr_3395 , wr_3391 , wr_3394 );
  not g3389( G330    ,           wr_2454 );
  nor g3390( wr_2435 , wr_2434 , wr_2432 );
  nor g3391( G321    , wr_2897 , wr_2895 );
  nor g3392( G338    , wr_3033 , wr_3031 );
  nor g3393( G370    , wr_3218 , wr_3216 );
  nor g3394( G399    , wr_3395 , wr_3393 );
  not g3395( G327    ,           wr_2435 );

endmodule
