// NOR_NOT mapped module c3540

module c3540 (
  input  G1      ,
  input  G13     ,
  input  G20     ,
  input  G33     ,
  input  G41     ,
  input  G45     ,
  input  G50     ,
  input  G58     ,
  input  G68     ,
  input  G77     ,
  input  G87     ,
  input  G97     ,
  input  G107    ,
  input  G116    ,
  input  G124    ,
  input  G125    ,
  input  G128    ,
  input  G132    ,
  input  G137    ,
  input  G143    ,
  input  G150    ,
  input  G159    ,
  input  G169    ,
  input  G179    ,
  input  G190    ,
  input  G200    ,
  input  G213    ,
  input  G222    ,
  input  G223    ,
  input  G226    ,
  input  G232    ,
  input  G238    ,
  input  G244    ,
  input  G250    ,
  input  G257    ,
  input  G264    ,
  input  G270    ,
  input  G274    ,
  input  G283    ,
  input  G294    ,
  input  G303    ,
  input  G311    ,
  input  G317    ,
  input  G322    ,
  input  G326    ,
  input  G329    ,
  input  G330    ,
  input  G343    ,
  input  G1698   ,
  input  G2897   ,
  output G353    ,
  output G355    ,
  output G361    ,
  output G358    ,
  output G351    ,
  output G372    ,
  output G369    ,
  output G399    ,
  output G364    ,
  output G396    ,
  output G384    ,
  output G367    ,
  output G387    ,
  output G393    ,
  output G390    ,
  output G378    ,
  output G375    ,
  output G381    ,
  output G407    ,
  output G409    ,
  output G405    ,
  output G402    );

  wire wr_23;
  wire wr_24;
  wire wr_25;
  wire wr_26;
  wire wr_27;
  wire wr_28;
  wire wr_29;
  wire wr_30;
  wire wr_31;
  wire wr_32;
  wire wr_33;
  wire wr_34;
  wire wr_35;
  wire wr_36;
  wire wr_37;
  wire wr_38;
  wire wr_39;
  wire wr_40;
  wire wr_41;
  wire wr_42;
  wire wr_43;
  wire wr_44;
  wire wr_45;
  wire wr_46;
  wire wr_47;
  wire wr_48;
  wire wr_49;
  wire wr_50;
  wire wr_51;
  wire wr_52;
  wire wr_53;
  wire wr_54;
  wire wr_55;
  wire wr_56;
  wire wr_57;
  wire wr_58;
  wire wr_59;
  wire wr_60;
  wire wr_61;
  wire wr_62;
  wire wr_63;
  wire wr_64;
  wire wr_65;
  wire wr_66;
  wire wr_67;
  wire wr_68;
  wire wr_69;
  wire wr_70;
  wire wr_71;
  wire wr_72;
  wire wr_73;
  wire wr_74;
  wire wr_75;
  wire wr_76;
  wire wr_77;
  wire wr_78;
  wire wr_79;
  wire wr_80;
  wire wr_81;
  wire wr_82;
  wire wr_83;
  wire wr_84;
  wire wr_85;
  wire wr_86;
  wire wr_87;
  wire wr_88;
  wire wr_89;
  wire wr_90;
  wire wr_91;
  wire wr_92;
  wire wr_93;
  wire wr_94;
  wire wr_95;
  wire wr_96;
  wire wr_97;
  wire wr_98;
  wire wr_99;
  wire wr_100;
  wire wr_101;
  wire wr_102;
  wire wr_103;
  wire wr_104;
  wire wr_105;
  wire wr_106;
  wire wr_107;
  wire wr_108;
  wire wr_109;
  wire wr_110;
  wire wr_111;
  wire wr_112;
  wire wr_113;
  wire wr_114;
  wire wr_115;
  wire wr_116;
  wire wr_117;
  wire wr_118;
  wire wr_119;
  wire wr_120;
  wire wr_121;
  wire wr_122;
  wire wr_123;
  wire wr_124;
  wire wr_125;
  wire wr_126;
  wire wr_127;
  wire wr_128;
  wire wr_129;
  wire wr_130;
  wire wr_131;
  wire wr_132;
  wire wr_133;
  wire wr_134;
  wire wr_135;
  wire wr_136;
  wire wr_137;
  wire wr_138;
  wire wr_139;
  wire wr_140;
  wire wr_141;
  wire wr_142;
  wire wr_143;
  wire wr_144;
  wire wr_145;
  wire wr_146;
  wire wr_147;
  wire wr_148;
  wire wr_149;
  wire wr_150;
  wire wr_151;
  wire wr_152;
  wire wr_153;
  wire wr_154;
  wire wr_155;
  wire wr_156;
  wire wr_157;
  wire wr_158;
  wire wr_159;
  wire wr_160;
  wire wr_161;
  wire wr_162;
  wire wr_163;
  wire wr_164;
  wire wr_165;
  wire wr_166;
  wire wr_167;
  wire wr_168;
  wire wr_169;
  wire wr_170;
  wire wr_171;
  wire wr_172;
  wire wr_173;
  wire wr_174;
  wire wr_175;
  wire wr_176;
  wire wr_177;
  wire wr_178;
  wire wr_179;
  wire wr_180;
  wire wr_181;
  wire wr_182;
  wire wr_183;
  wire wr_184;
  wire wr_185;
  wire wr_186;
  wire wr_187;
  wire wr_188;
  wire wr_189;
  wire wr_190;
  wire wr_191;
  wire wr_192;
  wire wr_193;
  wire wr_194;
  wire wr_195;
  wire wr_196;
  wire wr_197;
  wire wr_198;
  wire wr_199;
  wire wr_200;
  wire wr_201;
  wire wr_202;
  wire wr_203;
  wire wr_204;
  wire wr_205;
  wire wr_206;
  wire wr_207;
  wire wr_208;
  wire wr_209;
  wire wr_210;
  wire wr_211;
  wire wr_212;
  wire wr_213;
  wire wr_214;
  wire wr_215;
  wire wr_216;
  wire wr_217;
  wire wr_218;
  wire wr_219;
  wire wr_220;
  wire wr_221;
  wire wr_222;
  wire wr_223;
  wire wr_224;
  wire wr_225;
  wire wr_226;
  wire wr_227;
  wire wr_228;
  wire wr_229;
  wire wr_230;
  wire wr_231;
  wire wr_232;
  wire wr_233;
  wire wr_234;
  wire wr_235;
  wire wr_236;
  wire wr_237;
  wire wr_238;
  wire wr_239;
  wire wr_240;
  wire wr_241;
  wire wr_242;
  wire wr_243;
  wire wr_244;
  wire wr_245;
  wire wr_246;
  wire wr_247;
  wire wr_248;
  wire wr_249;
  wire wr_250;
  wire wr_251;
  wire wr_252;
  wire wr_253;
  wire wr_254;
  wire wr_255;
  wire wr_256;
  wire wr_257;
  wire wr_258;
  wire wr_259;
  wire wr_260;
  wire wr_261;
  wire wr_262;
  wire wr_263;
  wire wr_264;
  wire wr_265;
  wire wr_266;
  wire wr_267;
  wire wr_268;
  wire wr_269;
  wire wr_270;
  wire wr_271;
  wire wr_272;
  wire wr_273;
  wire wr_274;
  wire wr_275;
  wire wr_276;
  wire wr_277;
  wire wr_278;
  wire wr_279;
  wire wr_280;
  wire wr_281;
  wire wr_282;
  wire wr_283;
  wire wr_284;
  wire wr_285;
  wire wr_286;
  wire wr_287;
  wire wr_288;
  wire wr_289;
  wire wr_290;
  wire wr_291;
  wire wr_292;
  wire wr_293;
  wire wr_294;
  wire wr_295;
  wire wr_296;
  wire wr_297;
  wire wr_298;
  wire wr_299;
  wire wr_300;
  wire wr_301;
  wire wr_302;
  wire wr_303;
  wire wr_304;
  wire wr_305;
  wire wr_306;
  wire wr_307;
  wire wr_308;
  wire wr_309;
  wire wr_310;
  wire wr_311;
  wire wr_312;
  wire wr_313;
  wire wr_314;
  wire wr_315;
  wire wr_316;
  wire wr_317;
  wire wr_318;
  wire wr_319;
  wire wr_320;
  wire wr_321;
  wire wr_322;
  wire wr_323;
  wire wr_324;
  wire wr_325;
  wire wr_326;
  wire wr_327;
  wire wr_328;
  wire wr_329;
  wire wr_330;
  wire wr_331;
  wire wr_332;
  wire wr_333;
  wire wr_334;
  wire wr_335;
  wire wr_336;
  wire wr_337;
  wire wr_338;
  wire wr_339;
  wire wr_340;
  wire wr_341;
  wire wr_342;
  wire wr_343;
  wire wr_344;
  wire wr_345;
  wire wr_346;
  wire wr_347;
  wire wr_348;
  wire wr_349;
  wire wr_350;
  wire wr_351;
  wire wr_352;
  wire wr_353;
  wire wr_354;
  wire wr_355;
  wire wr_356;
  wire wr_357;
  wire wr_358;
  wire wr_359;
  wire wr_360;
  wire wr_361;
  wire wr_362;
  wire wr_363;
  wire wr_364;
  wire wr_365;
  wire wr_366;
  wire wr_367;
  wire wr_368;
  wire wr_369;
  wire wr_370;
  wire wr_371;
  wire wr_372;
  wire wr_373;
  wire wr_374;
  wire wr_375;
  wire wr_376;
  wire wr_377;
  wire wr_378;
  wire wr_379;
  wire wr_380;
  wire wr_381;
  wire wr_382;
  wire wr_383;
  wire wr_384;
  wire wr_385;
  wire wr_386;
  wire wr_387;
  wire wr_388;
  wire wr_389;
  wire wr_390;
  wire wr_391;
  wire wr_392;
  wire wr_393;
  wire wr_394;
  wire wr_395;
  wire wr_396;
  wire wr_397;
  wire wr_398;
  wire wr_399;
  wire wr_400;
  wire wr_401;
  wire wr_402;
  wire wr_403;
  wire wr_404;
  wire wr_405;
  wire wr_406;
  wire wr_407;
  wire wr_408;
  wire wr_409;
  wire wr_410;
  wire wr_411;
  wire wr_412;
  wire wr_413;
  wire wr_414;
  wire wr_415;
  wire wr_416;
  wire wr_417;
  wire wr_418;
  wire wr_419;
  wire wr_420;
  wire wr_421;
  wire wr_422;
  wire wr_423;
  wire wr_424;
  wire wr_425;
  wire wr_426;
  wire wr_427;
  wire wr_428;
  wire wr_429;
  wire wr_430;
  wire wr_431;
  wire wr_432;
  wire wr_433;
  wire wr_434;
  wire wr_435;
  wire wr_436;
  wire wr_437;
  wire wr_438;
  wire wr_439;
  wire wr_440;
  wire wr_441;
  wire wr_442;
  wire wr_443;
  wire wr_444;
  wire wr_445;
  wire wr_446;
  wire wr_447;
  wire wr_448;
  wire wr_449;
  wire wr_450;
  wire wr_451;
  wire wr_452;
  wire wr_453;
  wire wr_454;
  wire wr_455;
  wire wr_456;
  wire wr_457;
  wire wr_458;
  wire wr_459;
  wire wr_460;
  wire wr_461;
  wire wr_462;
  wire wr_463;
  wire wr_464;
  wire wr_465;
  wire wr_466;
  wire wr_467;
  wire wr_468;
  wire wr_469;
  wire wr_470;
  wire wr_471;
  wire wr_472;
  wire wr_473;
  wire wr_474;
  wire wr_475;
  wire wr_476;
  wire wr_477;
  wire wr_478;
  wire wr_479;
  wire wr_480;
  wire wr_481;
  wire wr_482;
  wire wr_483;
  wire wr_484;
  wire wr_485;
  wire wr_486;
  wire wr_487;
  wire wr_488;
  wire wr_489;
  wire wr_490;
  wire wr_491;
  wire wr_492;
  wire wr_493;
  wire wr_494;
  wire wr_495;
  wire wr_496;
  wire wr_497;
  wire wr_498;
  wire wr_499;
  wire wr_500;
  wire wr_501;
  wire wr_502;
  wire wr_503;
  wire wr_504;
  wire wr_505;
  wire wr_506;
  wire wr_507;
  wire wr_508;
  wire wr_509;
  wire wr_510;
  wire wr_511;
  wire wr_512;
  wire wr_513;
  wire wr_514;
  wire wr_515;
  wire wr_516;
  wire wr_517;
  wire wr_518;
  wire wr_519;
  wire wr_520;
  wire wr_521;
  wire wr_522;
  wire wr_523;
  wire wr_524;
  wire wr_525;
  wire wr_526;
  wire wr_527;
  wire wr_528;
  wire wr_529;
  wire wr_530;
  wire wr_531;
  wire wr_532;
  wire wr_533;
  wire wr_534;
  wire wr_535;
  wire wr_536;
  wire wr_537;
  wire wr_538;
  wire wr_539;
  wire wr_540;
  wire wr_541;
  wire wr_542;
  wire wr_543;
  wire wr_544;
  wire wr_545;
  wire wr_546;
  wire wr_547;
  wire wr_548;
  wire wr_549;
  wire wr_550;
  wire wr_551;
  wire wr_552;
  wire wr_553;
  wire wr_554;
  wire wr_555;
  wire wr_556;
  wire wr_557;
  wire wr_558;
  wire wr_559;
  wire wr_560;
  wire wr_561;
  wire wr_562;
  wire wr_563;
  wire wr_564;
  wire wr_565;
  wire wr_566;
  wire wr_567;
  wire wr_568;
  wire wr_569;
  wire wr_570;
  wire wr_571;
  wire wr_572;
  wire wr_573;
  wire wr_574;
  wire wr_575;
  wire wr_576;
  wire wr_577;
  wire wr_578;
  wire wr_579;
  wire wr_580;
  wire wr_581;
  wire wr_582;
  wire wr_583;
  wire wr_584;
  wire wr_585;
  wire wr_586;
  wire wr_587;
  wire wr_588;
  wire wr_589;
  wire wr_590;
  wire wr_591;
  wire wr_592;
  wire wr_593;
  wire wr_594;
  wire wr_595;
  wire wr_596;
  wire wr_597;
  wire wr_598;
  wire wr_599;
  wire wr_600;
  wire wr_601;
  wire wr_602;
  wire wr_603;
  wire wr_604;
  wire wr_605;
  wire wr_606;
  wire wr_607;
  wire wr_608;
  wire wr_609;
  wire wr_610;
  wire wr_611;
  wire wr_612;
  wire wr_613;
  wire wr_614;
  wire wr_615;
  wire wr_616;
  wire wr_617;
  wire wr_618;
  wire wr_619;
  wire wr_620;
  wire wr_621;
  wire wr_622;
  wire wr_623;
  wire wr_624;
  wire wr_625;
  wire wr_626;
  wire wr_627;
  wire wr_628;
  wire wr_629;
  wire wr_630;
  wire wr_631;
  wire wr_632;
  wire wr_633;
  wire wr_634;
  wire wr_635;
  wire wr_636;
  wire wr_637;
  wire wr_638;
  wire wr_639;
  wire wr_640;
  wire wr_641;
  wire wr_642;
  wire wr_643;
  wire wr_644;
  wire wr_645;
  wire wr_646;
  wire wr_647;
  wire wr_648;
  wire wr_649;
  wire wr_650;
  wire wr_651;
  wire wr_652;
  wire wr_653;
  wire wr_654;
  wire wr_655;
  wire wr_656;
  wire wr_657;
  wire wr_658;
  wire wr_659;
  wire wr_660;
  wire wr_661;
  wire wr_662;
  wire wr_663;
  wire wr_664;
  wire wr_665;
  wire wr_666;
  wire wr_667;
  wire wr_668;
  wire wr_669;
  wire wr_670;
  wire wr_671;
  wire wr_672;
  wire wr_673;
  wire wr_674;
  wire wr_675;
  wire wr_676;
  wire wr_677;
  wire wr_678;
  wire wr_679;
  wire wr_680;
  wire wr_681;
  wire wr_682;
  wire wr_683;
  wire wr_684;
  wire wr_685;
  wire wr_686;
  wire wr_687;
  wire wr_688;
  wire wr_689;
  wire wr_690;
  wire wr_691;
  wire wr_692;
  wire wr_693;
  wire wr_694;
  wire wr_695;
  wire wr_696;
  wire wr_697;
  wire wr_698;
  wire wr_699;
  wire wr_700;
  wire wr_701;
  wire wr_702;
  wire wr_703;
  wire wr_704;
  wire wr_705;
  wire wr_706;
  wire wr_707;
  wire wr_708;
  wire wr_709;
  wire wr_710;
  wire wr_711;
  wire wr_712;
  wire wr_713;
  wire wr_714;
  wire wr_715;
  wire wr_716;
  wire wr_717;
  wire wr_718;
  wire wr_719;
  wire wr_720;
  wire wr_721;
  wire wr_722;
  wire wr_723;
  wire wr_724;
  wire wr_725;
  wire wr_726;
  wire wr_727;
  wire wr_728;
  wire wr_729;
  wire wr_730;
  wire wr_731;
  wire wr_732;
  wire wr_733;
  wire wr_734;
  wire wr_735;
  wire wr_736;
  wire wr_737;
  wire wr_738;
  wire wr_739;
  wire wr_740;
  wire wr_741;
  wire wr_742;
  wire wr_743;
  wire wr_744;
  wire wr_745;
  wire wr_746;
  wire wr_747;
  wire wr_748;
  wire wr_749;
  wire wr_750;
  wire wr_751;
  wire wr_752;
  wire wr_753;
  wire wr_754;
  wire wr_755;
  wire wr_756;
  wire wr_757;
  wire wr_758;
  wire wr_759;
  wire wr_760;
  wire wr_761;
  wire wr_762;
  wire wr_763;
  wire wr_764;
  wire wr_765;
  wire wr_766;
  wire wr_767;
  wire wr_768;
  wire wr_769;
  wire wr_770;
  wire wr_771;
  wire wr_772;
  wire wr_773;
  wire wr_774;
  wire wr_775;
  wire wr_776;
  wire wr_777;
  wire wr_778;
  wire wr_779;
  wire wr_780;
  wire wr_781;
  wire wr_782;
  wire wr_783;
  wire wr_784;
  wire wr_785;
  wire wr_786;
  wire wr_787;
  wire wr_788;
  wire wr_789;
  wire wr_790;
  wire wr_791;
  wire wr_792;
  wire wr_793;
  wire wr_794;
  wire wr_795;
  wire wr_796;
  wire wr_797;
  wire wr_798;
  wire wr_799;
  wire wr_800;
  wire wr_801;
  wire wr_802;
  wire wr_803;
  wire wr_804;
  wire wr_805;
  wire wr_806;
  wire wr_807;
  wire wr_808;
  wire wr_809;
  wire wr_810;
  wire wr_811;
  wire wr_812;
  wire wr_813;
  wire wr_814;
  wire wr_815;
  wire wr_816;
  wire wr_817;
  wire wr_818;
  wire wr_819;
  wire wr_820;
  wire wr_821;
  wire wr_822;
  wire wr_823;
  wire wr_824;
  wire wr_825;
  wire wr_826;
  wire wr_827;
  wire wr_828;
  wire wr_829;
  wire wr_830;
  wire wr_831;
  wire wr_832;
  wire wr_833;
  wire wr_834;
  wire wr_835;
  wire wr_836;
  wire wr_837;
  wire wr_838;
  wire wr_839;
  wire wr_840;
  wire wr_841;
  wire wr_842;
  wire wr_843;
  wire wr_844;
  wire wr_845;
  wire wr_846;
  wire wr_847;
  wire wr_848;
  wire wr_849;
  wire wr_850;
  wire wr_851;
  wire wr_852;
  wire wr_853;
  wire wr_854;
  wire wr_855;
  wire wr_856;
  wire wr_857;
  wire wr_858;
  wire wr_859;
  wire wr_860;
  wire wr_861;
  wire wr_862;
  wire wr_863;
  wire wr_864;
  wire wr_865;
  wire wr_866;
  wire wr_867;
  wire wr_868;
  wire wr_869;
  wire wr_870;
  wire wr_871;
  wire wr_872;
  wire wr_873;
  wire wr_874;
  wire wr_875;
  wire wr_876;
  wire wr_877;
  wire wr_878;
  wire wr_879;
  wire wr_880;
  wire wr_881;
  wire wr_882;
  wire wr_883;
  wire wr_884;
  wire wr_885;
  wire wr_886;
  wire wr_887;
  wire wr_888;
  wire wr_889;
  wire wr_890;
  wire wr_891;
  wire wr_892;
  wire wr_893;
  wire wr_894;
  wire wr_895;
  wire wr_896;
  wire wr_897;
  wire wr_898;
  wire wr_899;
  wire wr_900;
  wire wr_901;
  wire wr_902;
  wire wr_903;
  wire wr_904;
  wire wr_905;
  wire wr_906;
  wire wr_907;
  wire wr_908;
  wire wr_909;
  wire wr_910;
  wire wr_911;
  wire wr_912;
  wire wr_913;
  wire wr_914;
  wire wr_915;
  wire wr_916;
  wire wr_917;
  wire wr_918;
  wire wr_919;
  wire wr_920;
  wire wr_921;
  wire wr_922;
  wire wr_923;
  wire wr_924;
  wire wr_925;
  wire wr_926;
  wire wr_927;
  wire wr_928;
  wire wr_929;
  wire wr_930;
  wire wr_931;
  wire wr_932;
  wire wr_933;
  wire wr_934;
  wire wr_935;
  wire wr_936;
  wire wr_937;
  wire wr_938;
  wire wr_939;
  wire wr_940;
  wire wr_941;
  wire wr_942;
  wire wr_943;
  wire wr_944;
  wire wr_945;
  wire wr_946;
  wire wr_947;
  wire wr_948;
  wire wr_949;
  wire wr_950;
  wire wr_951;
  wire wr_952;
  wire wr_953;
  wire wr_954;
  wire wr_955;
  wire wr_956;
  wire wr_957;
  wire wr_958;
  wire wr_959;
  wire wr_960;
  wire wr_961;
  wire wr_962;
  wire wr_963;
  wire wr_964;
  wire wr_965;
  wire wr_966;
  wire wr_967;
  wire wr_968;
  wire wr_969;
  wire wr_970;
  wire wr_971;
  wire wr_972;
  wire wr_973;
  wire wr_974;
  wire wr_975;
  wire wr_976;
  wire wr_977;
  wire wr_978;
  wire wr_979;
  wire wr_980;
  wire wr_981;
  wire wr_982;
  wire wr_983;
  wire wr_984;
  wire wr_985;
  wire wr_986;
  wire wr_987;
  wire wr_988;
  wire wr_989;
  wire wr_990;
  wire wr_991;
  wire wr_992;
  wire wr_993;
  wire wr_994;
  wire wr_995;
  wire wr_996;
  wire wr_997;
  wire wr_998;
  wire wr_999;
  wire wr_1000;
  wire wr_1001;
  wire wr_1002;
  wire wr_1003;
  wire wr_1004;
  wire wr_1005;
  wire wr_1006;
  wire wr_1007;
  wire wr_1008;
  wire wr_1009;
  wire wr_1010;
  wire wr_1011;
  wire wr_1012;
  wire wr_1013;
  wire wr_1014;
  wire wr_1015;
  wire wr_1016;
  wire wr_1017;
  wire wr_1018;
  wire wr_1019;
  wire wr_1020;
  wire wr_1021;
  wire wr_1022;
  wire wr_1023;
  wire wr_1024;
  wire wr_1025;
  wire wr_1026;
  wire wr_1027;
  wire wr_1028;
  wire wr_1029;
  wire wr_1030;
  wire wr_1031;
  wire wr_1032;
  wire wr_1033;
  wire wr_1034;
  wire wr_1035;
  wire wr_1036;
  wire wr_1037;
  wire wr_1038;
  wire wr_1039;
  wire wr_1040;
  wire wr_1041;
  wire wr_1042;
  wire wr_1043;
  wire wr_1044;
  wire wr_1045;
  wire wr_1046;
  wire wr_1047;
  wire wr_1048;
  wire wr_1049;
  wire wr_1050;
  wire wr_1051;
  wire wr_1052;
  wire wr_1053;
  wire wr_1054;
  wire wr_1055;
  wire wr_1056;
  wire wr_1057;
  wire wr_1058;
  wire wr_1059;
  wire wr_1060;
  wire wr_1061;
  wire wr_1062;
  wire wr_1063;
  wire wr_1064;
  wire wr_1065;
  wire wr_1066;
  wire wr_1067;
  wire wr_1068;
  wire wr_1069;
  wire wr_1070;
  wire wr_1071;
  wire wr_1072;
  wire wr_1073;
  wire wr_1074;
  wire wr_1075;
  wire wr_1076;
  wire wr_1077;
  wire wr_1078;
  wire wr_1079;
  wire wr_1080;
  wire wr_1081;
  wire wr_1082;
  wire wr_1083;
  wire wr_1084;
  wire wr_1085;
  wire wr_1086;
  wire wr_1087;
  wire wr_1088;
  wire wr_1089;
  wire wr_1090;
  wire wr_1091;
  wire wr_1092;
  wire wr_1093;
  wire wr_1094;
  wire wr_1095;
  wire wr_1096;
  wire wr_1097;
  wire wr_1098;
  wire wr_1099;
  wire wr_1100;
  wire wr_1101;
  wire wr_1102;
  wire wr_1103;
  wire wr_1104;
  wire wr_1105;
  wire wr_1106;
  wire wr_1107;
  wire wr_1108;
  wire wr_1109;
  wire wr_1110;
  wire wr_1111;
  wire wr_1112;
  wire wr_1113;
  wire wr_1114;
  wire wr_1115;
  wire wr_1116;
  wire wr_1117;
  wire wr_1118;
  wire wr_1119;
  wire wr_1120;
  wire wr_1121;
  wire wr_1122;
  wire wr_1123;
  wire wr_1124;
  wire wr_1125;
  wire wr_1126;
  wire wr_1127;
  wire wr_1128;
  wire wr_1129;
  wire wr_1130;
  wire wr_1131;
  wire wr_1132;
  wire wr_1133;
  wire wr_1134;
  wire wr_1135;
  wire wr_1136;
  wire wr_1137;
  wire wr_1138;
  wire wr_1139;
  wire wr_1140;
  wire wr_1141;
  wire wr_1142;
  wire wr_1143;
  wire wr_1144;
  wire wr_1145;
  wire wr_1146;
  wire wr_1147;
  wire wr_1148;
  wire wr_1149;
  wire wr_1150;
  wire wr_1151;
  wire wr_1152;
  wire wr_1153;
  wire wr_1154;
  wire wr_1155;
  wire wr_1156;
  wire wr_1157;
  wire wr_1158;
  wire wr_1159;
  wire wr_1160;
  wire wr_1161;
  wire wr_1162;
  wire wr_1163;
  wire wr_1164;
  wire wr_1165;
  wire wr_1166;
  wire wr_1167;
  wire wr_1168;
  wire wr_1169;
  wire wr_1170;
  wire wr_1171;
  wire wr_1172;
  wire wr_1173;
  wire wr_1174;
  wire wr_1175;
  wire wr_1176;
  wire wr_1177;
  wire wr_1178;
  wire wr_1179;
  wire wr_1180;
  wire wr_1181;
  wire wr_1182;
  wire wr_1183;
  wire wr_1184;
  wire wr_1185;
  wire wr_1186;
  wire wr_1187;
  wire wr_1188;
  wire wr_1189;
  wire wr_1190;
  wire wr_1191;
  wire wr_1192;
  wire wr_1193;
  wire wr_1194;
  wire wr_1195;
  wire wr_1196;
  wire wr_1197;
  wire wr_1198;
  wire wr_1199;
  wire wr_1200;
  wire wr_1201;
  wire wr_1202;
  wire wr_1203;
  wire wr_1204;
  wire wr_1205;
  wire wr_1206;
  wire wr_1207;
  wire wr_1208;
  wire wr_1209;
  wire wr_1210;
  wire wr_1211;
  wire wr_1212;
  wire wr_1213;
  wire wr_1214;
  wire wr_1215;
  wire wr_1216;
  wire wr_1217;
  wire wr_1218;
  wire wr_1219;
  wire wr_1220;
  wire wr_1221;
  wire wr_1222;
  wire wr_1223;
  wire wr_1224;
  wire wr_1225;
  wire wr_1226;
  wire wr_1227;
  wire wr_1228;
  wire wr_1229;
  wire wr_1230;
  wire wr_1231;
  wire wr_1232;
  wire wr_1233;
  wire wr_1234;
  wire wr_1235;
  wire wr_1236;
  wire wr_1237;
  wire wr_1238;
  wire wr_1239;
  wire wr_1240;
  wire wr_1241;
  wire wr_1242;
  wire wr_1243;
  wire wr_1244;
  wire wr_1245;
  wire wr_1246;
  wire wr_1247;
  wire wr_1248;
  wire wr_1249;
  wire wr_1250;
  wire wr_1251;
  wire wr_1252;
  wire wr_1253;
  wire wr_1254;
  wire wr_1255;
  wire wr_1256;
  wire wr_1257;
  wire wr_1258;
  wire wr_1259;
  wire wr_1260;
  wire wr_1261;
  wire wr_1262;
  wire wr_1263;
  wire wr_1264;
  wire wr_1265;
  wire wr_1266;
  wire wr_1267;
  wire wr_1268;
  wire wr_1269;
  wire wr_1270;
  wire wr_1271;
  wire wr_1272;
  wire wr_1273;
  wire wr_1274;
  wire wr_1275;
  wire wr_1276;
  wire wr_1277;
  wire wr_1278;
  wire wr_1279;
  wire wr_1280;
  wire wr_1281;
  wire wr_1282;
  wire wr_1283;
  wire wr_1284;
  wire wr_1285;
  wire wr_1286;
  wire wr_1287;
  wire wr_1288;
  wire wr_1289;
  wire wr_1290;
  wire wr_1291;
  wire wr_1292;
  wire wr_1293;
  wire wr_1294;
  wire wr_1295;
  wire wr_1296;
  wire wr_1297;
  wire wr_1298;
  wire wr_1299;
  wire wr_1300;
  wire wr_1301;
  wire wr_1302;
  wire wr_1303;
  wire wr_1304;
  wire wr_1305;
  wire wr_1306;
  wire wr_1307;
  wire wr_1308;
  wire wr_1309;
  wire wr_1310;
  wire wr_1311;
  wire wr_1312;
  wire wr_1313;
  wire wr_1314;
  wire wr_1315;
  wire wr_1316;
  wire wr_1317;
  wire wr_1318;
  wire wr_1319;
  wire wr_1320;
  wire wr_1321;
  wire wr_1322;
  wire wr_1323;
  wire wr_1324;
  wire wr_1325;
  wire wr_1326;
  wire wr_1327;
  wire wr_1328;
  wire wr_1329;
  wire wr_1330;
  wire wr_1331;
  wire wr_1332;
  wire wr_1333;
  wire wr_1334;
  wire wr_1335;
  wire wr_1336;
  wire wr_1337;
  wire wr_1338;
  wire wr_1339;
  wire wr_1340;
  wire wr_1341;
  wire wr_1342;
  wire wr_1343;
  wire wr_1344;
  wire wr_1345;
  wire wr_1346;
  wire wr_1347;
  wire wr_1348;
  wire wr_1349;
  wire wr_1350;
  wire wr_1351;
  wire wr_1352;
  wire wr_1353;
  wire wr_1354;
  wire wr_1355;
  wire wr_1356;
  wire wr_1357;
  wire wr_1358;
  wire wr_1359;
  wire wr_1360;
  wire wr_1361;
  wire wr_1362;
  wire wr_1363;
  wire wr_1364;
  wire wr_1365;
  wire wr_1366;
  wire wr_1367;
  wire wr_1368;
  wire wr_1369;
  wire wr_1370;
  wire wr_1371;
  wire wr_1372;
  wire wr_1373;
  wire wr_1374;
  wire wr_1375;
  wire wr_1376;
  wire wr_1377;
  wire wr_1378;
  wire wr_1379;
  wire wr_1380;
  wire wr_1381;
  wire wr_1382;
  wire wr_1383;
  wire wr_1384;
  wire wr_1385;
  wire wr_1386;
  wire wr_1387;
  wire wr_1388;
  wire wr_1389;
  wire wr_1390;
  wire wr_1391;
  wire wr_1392;
  wire wr_1393;
  wire wr_1394;
  wire wr_1395;
  wire wr_1396;
  wire wr_1397;
  wire wr_1398;
  wire wr_1399;
  wire wr_1400;
  wire wr_1401;
  wire wr_1402;
  wire wr_1403;
  wire wr_1404;
  wire wr_1405;
  wire wr_1406;
  wire wr_1407;
  wire wr_1408;
  wire wr_1409;
  wire wr_1410;
  wire wr_1411;
  wire wr_1412;
  wire wr_1413;
  wire wr_1414;
  wire wr_1415;
  wire wr_1416;
  wire wr_1417;
  wire wr_1418;
  wire wr_1419;
  wire wr_1420;
  wire wr_1421;
  wire wr_1422;
  wire wr_1423;
  wire wr_1424;
  wire wr_1425;
  wire wr_1426;
  wire wr_1427;
  wire wr_1428;
  wire wr_1429;
  wire wr_1430;
  wire wr_1431;
  wire wr_1432;
  wire wr_1433;
  wire wr_1434;
  wire wr_1435;
  wire wr_1436;
  wire wr_1437;
  wire wr_1438;
  wire wr_1439;
  wire wr_1440;
  wire wr_1441;
  wire wr_1442;
  wire wr_1443;
  wire wr_1444;
  wire wr_1445;
  wire wr_1446;
  wire wr_1447;
  wire wr_1448;
  wire wr_1449;
  wire wr_1450;
  wire wr_1451;
  wire wr_1452;
  wire wr_1453;
  wire wr_1454;
  wire wr_1455;
  wire wr_1456;
  wire wr_1457;
  wire wr_1458;
  wire wr_1459;
  wire wr_1460;
  wire wr_1461;
  wire wr_1462;
  wire wr_1463;
  wire wr_1464;
  wire wr_1465;
  wire wr_1466;
  wire wr_1467;
  wire wr_1468;
  wire wr_1469;
  wire wr_1470;
  wire wr_1471;
  wire wr_1472;
  wire wr_1473;
  wire wr_1474;
  wire wr_1475;
  wire wr_1476;
  wire wr_1477;
  wire wr_1478;
  wire wr_1479;
  wire wr_1480;
  wire wr_1481;
  wire wr_1482;
  wire wr_1483;
  wire wr_1484;
  wire wr_1485;
  wire wr_1486;
  wire wr_1487;
  wire wr_1488;
  wire wr_1489;
  wire wr_1490;
  wire wr_1491;
  wire wr_1492;
  wire wr_1493;
  wire wr_1494;
  wire wr_1495;
  wire wr_1496;
  wire wr_1497;
  wire wr_1498;
  wire wr_1499;
  wire wr_1500;
  wire wr_1501;
  wire wr_1502;
  wire wr_1503;
  wire wr_1504;
  wire wr_1505;
  wire wr_1506;
  wire wr_1507;
  wire wr_1508;
  wire wr_1509;
  wire wr_1510;
  wire wr_1511;
  wire wr_1512;
  wire wr_1513;
  wire wr_1514;
  wire wr_1515;
  wire wr_1516;
  wire wr_1517;
  wire wr_1518;
  wire wr_1519;
  wire wr_1520;
  wire wr_1521;
  wire wr_1522;
  wire wr_1523;
  wire wr_1524;
  wire wr_1525;
  wire wr_1526;
  wire wr_1527;
  wire wr_1528;
  wire wr_1529;
  wire wr_1530;
  wire wr_1531;
  wire wr_1532;
  wire wr_1533;
  wire wr_1534;
  wire wr_1535;
  wire wr_1536;
  wire wr_1537;
  wire wr_1538;
  wire wr_1539;
  wire wr_1540;
  wire wr_1541;
  wire wr_1542;
  wire wr_1543;
  wire wr_1544;
  wire wr_1545;
  wire wr_1546;
  wire wr_1547;
  wire wr_1548;
  wire wr_1549;
  wire wr_1550;
  wire wr_1551;
  wire wr_1552;
  wire wr_1553;
  wire wr_1554;
  wire wr_1555;
  wire wr_1556;
  wire wr_1557;
  wire wr_1558;
  wire wr_1559;
  wire wr_1560;
  wire wr_1561;
  wire wr_1562;
  wire wr_1563;
  wire wr_1564;
  wire wr_1565;
  wire wr_1566;
  wire wr_1567;
  wire wr_1568;
  wire wr_1569;
  wire wr_1570;
  wire wr_1571;
  wire wr_1572;
  wire wr_1573;
  wire wr_1574;
  wire wr_1575;
  wire wr_1576;
  wire wr_1577;
  wire wr_1578;
  wire wr_1579;
  wire wr_1580;

  nor    g1( wr_23   , G68     , G50     );
  not    g2( wr_27   ,           G87     );
  not    g3( wr_30   ,           G1      );
  not    g4( wr_31   ,           G20     );
  not    g5( wr_36   ,           G250    );
  not    g6( wr_41   ,           G58     );
  not    g7( wr_42   ,           G232    );
  not    g8( wr_44   ,           G50     );
  not    g9( wr_45   ,           G226    );
  not   g10( wr_47   ,           G77     );
  not   g11( wr_48   ,           G244    );
  not   g12( wr_50   ,           G68     );
  not   g13( wr_51   ,           G238    );
  not   g14( wr_59   ,           G97     );
  not   g15( wr_60   ,           G257    );
  not   g16( wr_63   ,           G116    );
  not   g17( wr_64   ,           G270    );
  not   g18( wr_66   ,           G107    );
  not   g19( wr_67   ,           G264    );
  not   g20( wr_76   ,           G13     );
  not   g21( wr_146  ,           G33     );
  nor   g22( wr_162  , G33     , G20     );
  not   g23( wr_177  ,           G169    );
  not   g24( wr_178  ,           G274    );
  not   g25( wr_179  ,           G41     );
  not   g26( wr_184  ,           G45     );
  nor   g27( wr_185  , G41     , G1      );
  nor   g28( wr_193  , G1698   , G33     );
  not   g29( wr_199  ,           G283    );
  not   g30( wr_214  ,           G179    );
  not   g31( wr_222  ,           G200    );
  not   g32( wr_226  ,           G190    );
  nor   g33( wr_239  , G107    , G87     );
  not   g34( wr_303  ,           G303    );
  not   g35( wr_348  ,           G294    );
  not   g36( wr_389  ,           G159    );
  nor   g37( wr_403  , G45     , G41     );
  not   g38( wr_409  ,           G223    );
  not   g39( wr_447  ,           G150    );
  not   g40( wr_457  ,           G222    );
  not   g41( wr_613  ,           G213    );
  not   g42( wr_614  ,           G343    );
  nor   g43( wr_615  , G20     , G1      );
  not   g44( wr_1296 ,           G125    );
  not   g45( wr_1302 ,           G128    );
  not   g46( wr_839  ,           G132    );
  not   g47( wr_845  ,           G137    );
  not   g48( wr_847  ,           G143    );
  not   g49( wr_776  ,           G311    );
  not   g50( wr_778  ,           G317    );
  not   g51( wr_780  ,           G326    );
  not   g52( wr_782  ,           G322    );
  not   g53( wr_1405 ,           G124    );
  nor   g54( wr_128  , G58     , G50     );
  nor   g55( wr_1399 , G41     , G33     );
  nor   g56( wr_82   , G68     , G58     );
  not   g57( wr_641  ,           G330    );
  nor   g58( wr_689  , G33     , G13     );
  not   g59( wr_772  ,           G329    );
  nor   g60( wr_28   , G107    , G97     );
  not   g61( wr_1543 ,           G2897   );
  nor   g62( wr_37   , G264    , G257    );
  not   g63( wr_24   ,           wr_23   );
  nor   g64( wr_141  , wr_31   , wr_76   );
  nor   g65( wr_147  , wr_146  , G1      );
  nor   g66( wr_148  , wr_76   , wr_30   );
  nor   g67( wr_149  , wr_146  , wr_30   );
  nor   g68( wr_159  , wr_146  , G20     );
  not   g69( wr_163  ,           wr_162  );
  nor   g70( wr_165  , wr_66   , G97     );
  nor   g71( wr_166  , G107    , wr_59   );
  nor   g72( wr_180  , wr_179  , wr_146  );
  not   g73( wr_186  ,           wr_185  );
  not   g74( wr_194  ,           wr_193  );
  nor   g75( wr_196  , wr_193  , G33     );
  nor   g76( wr_200  , wr_199  , wr_146  );
  not   g77( wr_240  ,           wr_239  );
  nor   g78( wr_250  , wr_184  , G1      );
  nor   g79( wr_257  , wr_63   , wr_146  );
  nor   g80( wr_293  , wr_63   , wr_31   );
  nor   g81( wr_304  , wr_303  , wr_146  );
  nor   g82( wr_338  , G107    , wr_31   );
  nor   g83( wr_349  , wr_348  , wr_146  );
  nor   g84( wr_384  , wr_31   , G1      );
  nor   g85( wr_391  , wr_50   , G58     );
  nor   g86( wr_392  , G68     , wr_41   );
  nor   g87( wr_404  , wr_403  , G1      );
  nor   g88( wr_412  , wr_27   , wr_146  );
  nor   g89( wr_460  , wr_47   , wr_146  );
  nor   g90( wr_494  , wr_47   , wr_31   );
  nor   g91( wr_504  , wr_66   , wr_146  );
  nor   g92( wr_538  , G68     , wr_31   );
  nor   g93( wr_548  , wr_59   , wr_146  );
  not   g94( wr_616  ,           wr_615  );
  nor   g95( wr_718  , G190    , wr_31   );
  nor   g96( wr_720  , wr_214  , wr_31   );
  nor   g97( wr_721  , wr_222  , wr_31   );
  nor   g98( wr_32   , wr_31   , wr_30   );
  nor   g99( wr_99   , wr_48   , G238    );
  nor  g100( wr_100  , G244    , wr_51   );
  nor  g101( wr_102  , wr_42   , G226    );
  nor  g102( wr_103  , G232    , wr_45   );
  nor  g103( wr_1107 , wr_41   , G50     );
  nor  g104( wr_125  , G77     , wr_50   );
  nor  g105( wr_126  , wr_47   , G68     );
  nor  g106( wr_129  , wr_41   , wr_44   );
  nor  g107( wr_710  , G169    , wr_31   );
  nor  g108( wr_1376 , G41     , wr_146  );
  nor  g109( wr_88   , wr_64   , G264    );
  nor  g110( wr_89   , G270    , wr_67   );
  nor  g111( wr_91   , wr_60   , G250    );
  nor  g112( wr_92   , G257    , wr_36   );
  nor  g113( wr_114  , G116    , wr_66   );
  nor  g114( wr_115  , wr_63   , G107    );
  nor  g115( wr_117  , G97     , wr_27   );
  nor  g116( wr_118  , wr_59   , G87     );
  nor  g117( wr_1106 , wr_47   , wr_50   );
  not  g118( wr_1403 ,           wr_1399 );
  nor  g119( wr_83   , wr_82   , wr_44   );
  nor  g120( wr_671  , G41     , wr_31   );
  nor  g121( wr_805  , wr_184  , wr_76   );
  not  g122( wr_690  ,           wr_689  );
  nor  g123( wr_29   , wr_28   , wr_27   );
  nor  g124( wr_1515 , G343    , wr_613  );
  nor  g125( wr_49   , wr_48   , wr_47   );
  nor  g126( wr_52   , wr_51   , wr_50   );
  nor  g127( wr_65   , wr_64   , wr_63   );
  nor  g128( wr_68   , wr_67   , wr_66   );
  nor  g129( wr_46   , wr_45   , wr_44   );
  nor  g130( wr_62   , wr_36   , wr_27   );
  nor  g131( wr_43   , wr_42   , wr_41   );
  nor  g132( wr_61   , wr_60   , wr_59   );
  nor  g133( wr_955  , G13     , wr_30   );
  nor  g134( wr_963  , wr_50   , G50     );
  nor  g135( wr_38   , wr_37   , wr_36   );
  nor  g136( wr_25   , wr_24   , G58     );
  not  g137( wr_142  ,           wr_141  );
  not  g138( wr_150  ,           wr_149  );
  not  g139( wr_160  ,           wr_159  );
  nor  g140( wr_164  , wr_163  , wr_47   );
  nor  g141( wr_167  , wr_166  , wr_165  );
  nor  g142( wr_181  , wr_180  , wr_30   );
  nor  g143( wr_187  , wr_186  , wr_184  );
  nor  g144( wr_195  , wr_194  , wr_48   );
  not  g145( wr_197  ,           wr_196  );
  nor  g146( wr_238  , wr_163  , wr_50   );
  nor  g147( wr_241  , wr_240  , G97     );
  not  g148( wr_251  ,           wr_250  );
  nor  g149( wr_255  , wr_194  , wr_51   );
  nor  g150( wr_292  , wr_163  , wr_59   );
  nor  g151( wr_301  , wr_194  , wr_60   );
  nor  g152( wr_337  , wr_163  , wr_27   );
  nor  g153( wr_346  , wr_194  , wr_36   );
  nor  g154( wr_390  , wr_163  , wr_389  );
  nor  g155( wr_393  , wr_392  , wr_391  );
  not  g156( wr_405  ,           wr_404  );
  nor  g157( wr_410  , wr_194  , wr_409  );
  nor  g158( wr_448  , wr_163  , wr_447  );
  nor  g159( wr_458  , wr_194  , wr_457  );
  nor  g160( wr_493  , wr_163  , wr_41   );
  nor  g161( wr_502  , wr_194  , wr_42   );
  nor  g162( wr_537  , wr_163  , wr_44   );
  nor  g163( wr_546  , wr_194  , wr_45   );
  nor  g164( wr_617  , wr_616  , wr_76   );
  not  g165( wr_719  ,           wr_718  );
  not  g166( wr_739  ,           wr_720  );
  not  g167( wr_722  ,           wr_721  );
  nor  g168( wr_728  , wr_721  , wr_720  );
  not  g169( wr_33   ,           wr_32   );
  nor  g170( wr_101  , wr_100  , wr_99   );
  nor  g171( wr_104  , wr_103  , wr_102  );
  not  g172( wr_1108 ,           wr_1107 );
  nor  g173( wr_127  , wr_126  , wr_125  );
  nor  g174( wr_130  , wr_129  , wr_128  );
  nor  g175( wr_711  , wr_710  , wr_30   );
  nor  g176( wr_1400 , wr_1399 , wr_1376 );
  nor  g177( wr_90   , wr_89   , wr_88   );
  nor  g178( wr_93   , wr_92   , wr_91   );
  nor  g179( wr_116  , wr_115  , wr_114  );
  nor  g180( wr_119  , wr_118  , wr_117  );
  not  g181( wr_84   ,           wr_83   );
  not  g182( wr_1377 ,           wr_1376 );
  not  g183( wr_672  ,           wr_671  );
  not  g184( wr_806  ,           wr_805  );
  nor  g185( wr_691  , wr_690  , G20     );
  not  g186( wr_1516 ,           wr_1515 );
  nor  g187( wr_53   , wr_52   , wr_49   );
  nor  g188( wr_69   , wr_68   , wr_65   );
  not  g189( wr_959  ,           wr_955  );
  not  g190( wr_39   ,           wr_38   );
  not  g191( G355    ,           wr_29   );
  nor  g192( wr_143  , wr_142  , G1      );
  nor  g193( wr_151  , wr_150  , wr_31   );
  nor  g194( wr_161  , wr_160  , wr_66   );
  not  g195( wr_168  ,           wr_167  );
  not  g196( wr_182  ,           wr_181  );
  not  g197( wr_188  ,           wr_187  );
  nor  g198( wr_198  , wr_197  , wr_36   );
  nor  g199( wr_237  , wr_160  , wr_59   );
  nor  g200( wr_242  , wr_241  , wr_31   );
  nor  g201( wr_256  , wr_197  , wr_48   );
  nor  g202( wr_291  , wr_160  , wr_199  );
  nor  g203( wr_294  , wr_293  , wr_292  );
  nor  g204( wr_302  , wr_197  , wr_67   );
  nor  g205( wr_336  , wr_160  , wr_63   );
  nor  g206( wr_339  , wr_338  , wr_337  );
  nor  g207( wr_347  , wr_197  , wr_60   );
  nor  g208( wr_388  , wr_160  , wr_50   );
  not  g209( wr_394  ,           wr_393  );
  nor  g210( wr_411  , wr_197  , wr_45   );
  nor  g211( wr_446  , wr_160  , wr_41   );
  nor  g212( wr_449  , wr_25   , wr_31   );
  nor  g213( wr_459  , wr_197  , wr_409  );
  nor  g214( wr_492  , wr_160  , wr_27   );
  nor  g215( wr_495  , wr_494  , wr_493  );
  nor  g216( wr_503  , wr_197  , wr_51   );
  nor  g217( wr_536  , wr_160  , wr_47   );
  nor  g218( wr_539  , wr_538  , wr_537  );
  nor  g219( wr_547  , wr_197  , wr_42   );
  not  g220( wr_618  ,           wr_617  );
  nor  g221( wr_740  , wr_739  , G200    );
  nor  g222( wr_745  , wr_739  , wr_222  );
  nor  g223( wr_723  , wr_722  , wr_720  );
  not  g224( wr_729  ,           wr_728  );
  not  g225( wr_668  ,           wr_241  );
  nor  g226( wr_34   , wr_33   , G13     );
  not  g227( wr_105  ,           wr_104  );
  not  g228( wr_107  ,           wr_101  );
  not  g229( wr_131  ,           wr_130  );
  not  g230( wr_133  ,           wr_127  );
  not  g231( wr_712  ,           wr_711  );
  not  g232( wr_1401 ,           wr_1400 );
  not  g233( wr_94   ,           wr_93   );
  not  g234( wr_96   ,           wr_90   );
  not  g235( wr_120  ,           wr_119  );
  not  g236( wr_122  ,           wr_116  );
  nor  g237( wr_703  , wr_84   , G45     );
  nor  g238( wr_673  , wr_672  , wr_30   );
  nor  g239( wr_807  , wr_806  , G20     );
  not  g240( wr_692  ,           wr_691  );
  nor  g241( wr_1544 , wr_1516 , wr_1543 );
  not  g242( wr_54   ,           wr_53   );
  not  g243( wr_70   ,           wr_69   );
  nor  g244( wr_960  , wr_393  , wr_44   );
  nor  g245( wr_77   , wr_33   , wr_76   );
  nor  g246( wr_897  , wr_167  , wr_63   );
  not  g247( wr_26   ,           wr_25   );
  not  g248( wr_144  ,           wr_143  );
  nor  g249( wr_152  , wr_151  , wr_148  );
  nor  g250( wr_169  , wr_168  , wr_31   );
  nor  g251( wr_183  , wr_182  , wr_76   );
  nor  g252( wr_201  , wr_200  , wr_198  );
  nor  g253( wr_243  , wr_242  , wr_238  );
  nor  g254( wr_258  , wr_257  , wr_256  );
  not  g255( wr_295  ,           wr_294  );
  nor  g256( wr_305  , wr_304  , wr_302  );
  not  g257( wr_340  ,           wr_339  );
  nor  g258( wr_350  , wr_349  , wr_347  );
  nor  g259( wr_395  , wr_394  , wr_31   );
  nor  g260( wr_413  , wr_412  , wr_411  );
  nor  g261( wr_450  , wr_449  , wr_448  );
  nor  g262( wr_461  , wr_460  , wr_459  );
  not  g263( wr_496  ,           wr_495  );
  nor  g264( wr_505  , wr_504  , wr_503  );
  not  g265( wr_540  ,           wr_539  );
  nor  g266( wr_549  , wr_548  , wr_547  );
  nor  g267( wr_619  , wr_618  , wr_614  );
  not  g268( wr_741  ,           wr_740  );
  not  g269( wr_746  ,           wr_745  );
  nor  g270( wr_900  , wr_618  , wr_613  );
  not  g271( wr_724  ,           wr_723  );
  nor  g272( wr_733  , wr_729  , wr_718  );
  nor  g273( wr_730  , wr_729  , wr_719  );
  nor  g274( wr_669  , wr_668  , G116    );
  not  g275( wr_35   ,           wr_34   );
  nor  g276( wr_106  , wr_105  , wr_101  );
  nor  g277( wr_108  , wr_104  , wr_107  );
  nor  g278( wr_132  , wr_131  , wr_127  );
  nor  g279( wr_134  , wr_130  , wr_133  );
  nor  g280( wr_713  , wr_712  , wr_76   );
  nor  g281( wr_1402 , wr_1401 , G50     );
  nor  g282( wr_95   , wr_94   , wr_90   );
  nor  g283( wr_97   , wr_93   , wr_96   );
  nor  g284( wr_121  , wr_120  , wr_116  );
  nor  g285( wr_123  , wr_119  , wr_122  );
  not  g286( wr_674  ,           wr_673  );
  nor  g287( wr_808  , wr_807  , wr_30   );
  not  g288( wr_1551 ,           wr_1544 );
  nor  g289( wr_55   , wr_54   , wr_46   );
  nor  g290( wr_71   , wr_70   , wr_62   );
  not  g291( wr_961  ,           wr_960  );
  nor  g292( wr_956  , wr_955  , wr_77   );
  nor  g293( wr_78   , wr_77   , wr_34   );
  not  g294( wr_81   ,           wr_77   );
  not  g295( wr_898  ,           wr_897  );
  nor  g296( G353    , wr_26   , G77     );
  nor  g297( wr_145  , wr_144  , G97     );
  not  g298( wr_153  ,           wr_152  );
  nor  g299( wr_170  , wr_169  , wr_164  );
  nor  g300( wr_189  , wr_188  , wr_183  );
  not  g301( wr_192  ,           wr_183  );
  not  g302( wr_202  ,           wr_201  );
  nor  g303( wr_205  , wr_187  , wr_183  );
  nor  g304( wr_233  , wr_144  , G87     );
  not  g305( wr_244  ,           wr_243  );
  nor  g306( wr_252  , wr_251  , wr_183  );
  not  g307( wr_259  ,           wr_258  );
  nor  g308( wr_262  , wr_250  , wr_183  );
  nor  g309( wr_287  , wr_144  , G116    );
  nor  g310( wr_296  , wr_295  , wr_291  );
  not  g311( wr_306  ,           wr_305  );
  nor  g312( wr_332  , wr_144  , G107    );
  nor  g313( wr_341  , wr_340  , wr_336  );
  not  g314( wr_351  ,           wr_350  );
  nor  g315( wr_383  , wr_144  , G58     );
  nor  g316( wr_396  , wr_395  , wr_390  );
  nor  g317( wr_406  , wr_405  , wr_183  );
  not  g318( wr_414  ,           wr_413  );
  nor  g319( wr_417  , wr_404  , wr_183  );
  nor  g320( wr_442  , wr_144  , G50     );
  not  g321( wr_451  ,           wr_450  );
  not  g322( wr_462  ,           wr_461  );
  nor  g323( wr_488  , wr_144  , G77     );
  nor  g324( wr_497  , wr_496  , wr_492  );
  not  g325( wr_506  ,           wr_505  );
  nor  g326( wr_532  , wr_144  , G68     );
  nor  g327( wr_541  , wr_540  , wr_536  );
  not  g328( wr_550  ,           wr_549  );
  not  g329( wr_620  ,           wr_619  );
  nor  g330( wr_750  , wr_746  , wr_718  );
  nor  g331( wr_753  , wr_741  , wr_718  );
  nor  g332( wr_747  , wr_746  , wr_719  );
  not  g333( wr_901  ,           wr_900  );
  nor  g334( wr_742  , wr_741  , wr_719  );
  nor  g335( wr_736  , wr_724  , wr_718  );
  not  g336( wr_734  ,           wr_733  );
  not  g337( wr_731  ,           wr_730  );
  nor  g338( wr_725  , wr_724  , wr_719  );
  not  g339( wr_670  ,           wr_669  );
  nor  g340( wr_109  , wr_108  , wr_106  );
  nor  g341( wr_694  , wr_35   , G33     );
  nor  g342( wr_697  , wr_35   , wr_146  );
  nor  g343( wr_135  , wr_134  , wr_132  );
  nor  g344( wr_835  , wr_713  , wr_689  );
  nor  g345( wr_98   , wr_97   , wr_95   );
  nor  g346( wr_124  , wr_123  , wr_121  );
  not  g347( wr_717  ,           wr_713  );
  nor  g348( wr_675  , wr_674  , G13     );
  nor  g349( wr_714  , wr_713  , wr_691  );
  not  g350( wr_809  ,           wr_808  );
  not  g351( wr_56   ,           wr_55   );
  not  g352( wr_72   ,           wr_71   );
  nor  g353( wr_962  , wr_961  , wr_47   );
  not  g354( wr_957  ,           wr_956  );
  not  g355( wr_79   ,           wr_78   );
  nor  g356( wr_85   , wr_84   , wr_81   );
  nor  g357( wr_899  , wr_898  , wr_81   );
  nor  g358( wr_40   , wr_39   , wr_35   );
  nor  g359( wr_154  , wr_153  , wr_143  );
  not  g360( wr_171  ,           wr_170  );
  not  g361( wr_190  ,           wr_189  );
  nor  g362( wr_203  , wr_202  , wr_195  );
  not  g363( wr_206  ,           wr_205  );
  nor  g364( wr_245  , wr_244  , wr_237  );
  not  g365( wr_253  ,           wr_252  );
  nor  g366( wr_260  , wr_259  , wr_255  );
  not  g367( wr_263  ,           wr_262  );
  nor  g368( wr_297  , wr_296  , wr_152  );
  nor  g369( wr_307  , wr_306  , wr_301  );
  nor  g370( wr_342  , wr_341  , wr_152  );
  nor  g371( wr_352  , wr_351  , wr_346  );
  not  g372( wr_397  ,           wr_396  );
  not  g373( wr_407  ,           wr_406  );
  nor  g374( wr_415  , wr_414  , wr_410  );
  not  g375( wr_418  ,           wr_417  );
  nor  g376( wr_452  , wr_451  , wr_446  );
  nor  g377( wr_463  , wr_462  , wr_458  );
  nor  g378( wr_498  , wr_497  , wr_152  );
  nor  g379( wr_507  , wr_506  , wr_502  );
  nor  g380( wr_542  , wr_541  , wr_152  );
  nor  g381( wr_551  , wr_550  , wr_546  );
  nor  g382( wr_621  , wr_620  , wr_613  );
  not  g383( wr_751  ,           wr_750  );
  not  g384( wr_754  ,           wr_753  );
  not  g385( wr_748  ,           wr_747  );
  not  g386( wr_743  ,           wr_742  );
  not  g387( wr_737  ,           wr_736  );
  nor  g388( wr_1407 , wr_734  , wr_447  );
  nor  g389( wr_735  , wr_734  , wr_59   );
  nor  g390( wr_841  , wr_734  , wr_41   );
  nor  g391( wr_1122 , wr_734  , wr_27   );
  nor  g392( wr_1449 , wr_734  , wr_44   );
  nor  g393( wr_1041 , wr_734  , wr_50   );
  nor  g394( wr_1191 , wr_734  , wr_47   );
  nor  g395( wr_1298 , wr_734  , wr_389  );
  nor  g396( wr_1406 , wr_731  , wr_1405 );
  not  g397( wr_726  ,           wr_725  );
  nor  g398( wr_840  , wr_731  , wr_839  );
  nor  g399( wr_865  , wr_731  , wr_776  );
  nor  g400( wr_1448 , wr_731  , wr_1302 );
  nor  g401( wr_1470 , wr_731  , wr_303  );
  nor  g402( wr_1297 , wr_731  , wr_1296 );
  nor  g403( wr_1320 , wr_731  , wr_348  );
  nor  g404( wr_1379 , wr_731  , wr_199  );
  nor  g405( wr_1064 , wr_734  , wr_66   );
  nor  g406( wr_1109 , wr_1108 , wr_670  );
  nor  g407( wr_1213 , wr_734  , wr_63   );
  nor  g408( wr_774  , wr_734  , wr_348  );
  nor  g409( wr_1040 , wr_731  , wr_845  );
  nor  g410( wr_1063 , wr_731  , wr_778  );
  nor  g411( wr_1145 , wr_734  , wr_199  );
  nor  g412( wr_1190 , wr_731  , wr_847  );
  nor  g413( wr_1212 , wr_731  , wr_782  );
  not  g414( wr_110  ,           wr_109  );
  nor  g415( wr_698  , wr_697  , wr_694  );
  not  g416( wr_701  ,           wr_697  );
  nor  g417( wr_702  , wr_135  , wr_184  );
  nor  g418( wr_732  , wr_731  , wr_389  );
  nor  g419( wr_773  , wr_731  , wr_772  );
  not  g420( wr_836  ,           wr_835  );
  nor  g421( wr_1121 , wr_731  , wr_447  );
  nor  g422( wr_1144 , wr_731  , wr_780  );
  not  g423( wr_695  ,           wr_694  );
  not  g424( wr_715  ,           wr_714  );
  nor  g425( wr_810  , wr_809  , wr_675  );
  not  g426( wr_679  ,           wr_675  );
  nor  g427( wr_57   , wr_56   , wr_43   );
  nor  g428( wr_73   , wr_72   , wr_61   );
  nor  g429( wr_676  , wr_675  , wr_30   );
  nor  g430( wr_964  , wr_963  , wr_962  );
  not  g431( wr_136  ,           wr_135  );
  not  g432( wr_138  ,           wr_124  );
  not  g433( wr_112  ,           wr_98   );
  not  g434( wr_155  ,           wr_154  );
  nor  g435( wr_172  , wr_171  , wr_161  );
  nor  g436( wr_191  , wr_190  , wr_178  );
  nor  g437( wr_204  , wr_203  , wr_192  );
  nor  g438( wr_207  , wr_206  , wr_60   );
  nor  g439( wr_246  , wr_245  , wr_152  );
  nor  g440( wr_254  , wr_253  , wr_178  );
  nor  g441( wr_261  , wr_260  , wr_192  );
  nor  g442( wr_264  , wr_263  , wr_36   );
  nor  g443( wr_308  , wr_307  , wr_192  );
  nor  g444( wr_309  , wr_206  , wr_64   );
  nor  g445( wr_353  , wr_352  , wr_192  );
  nor  g446( wr_354  , wr_206  , wr_67   );
  nor  g447( wr_398  , wr_397  , wr_388  );
  nor  g448( wr_408  , wr_407  , wr_178  );
  nor  g449( wr_416  , wr_415  , wr_192  );
  nor  g450( wr_419  , wr_418  , wr_42   );
  nor  g451( wr_453  , wr_452  , wr_152  );
  nor  g452( wr_464  , wr_463  , wr_192  );
  nor  g453( wr_465  , wr_418  , wr_45   );
  nor  g454( wr_508  , wr_507  , wr_192  );
  nor  g455( wr_509  , wr_418  , wr_48   );
  nor  g456( wr_552  , wr_551  , wr_192  );
  nor  g457( wr_553  , wr_418  , wr_51   );
  not  g458( wr_623  ,           wr_621  );
  nor  g459( wr_1411 , wr_751  , wr_1296 );
  nor  g460( wr_1412 , wr_754  , wr_1302 );
  nor  g461( wr_846  , wr_751  , wr_845  );
  nor  g462( wr_848  , wr_754  , wr_847  );
  nor  g463( wr_869  , wr_751  , wr_303  );
  nor  g464( wr_870  , wr_754  , wr_348  );
  nor  g465( wr_1453 , wr_751  , wr_839  );
  nor  g466( wr_1454 , wr_754  , wr_845  );
  nor  g467( wr_1474 , wr_751  , wr_348  );
  nor  g468( wr_1475 , wr_754  , wr_199  );
  nor  g469( wr_1303 , wr_751  , wr_1302 );
  nor  g470( wr_1304 , wr_754  , wr_839  );
  nor  g471( wr_1323 , wr_751  , wr_199  );
  nor  g472( wr_1324 , wr_754  , wr_63   );
  nor  g473( wr_1382 , wr_751  , wr_63   );
  nor  g474( wr_1383 , wr_754  , wr_66   );
  nor  g475( wr_1410 , wr_748  , wr_839  );
  nor  g476( wr_844  , wr_748  , wr_447  );
  nor  g477( wr_868  , wr_748  , wr_199  );
  nor  g478( wr_1452 , wr_748  , wr_847  );
  nor  g479( wr_1473 , wr_748  , wr_63   );
  nor  g480( wr_1301 , wr_748  , wr_845  );
  nor  g481( wr_1322 , wr_748  , wr_66   );
  nor  g482( wr_1381 , wr_748  , wr_59   );
  nor  g483( wr_1409 , wr_743  , wr_845  );
  nor  g484( wr_843  , wr_743  , wr_389  );
  nor  g485( wr_867  , wr_743  , wr_63   );
  nor  g486( wr_1045 , wr_751  , wr_847  );
  nor  g487( wr_1046 , wr_754  , wr_447  );
  nor  g488( wr_1068 , wr_751  , wr_776  );
  nor  g489( wr_1069 , wr_754  , wr_303  );
  nor  g490( wr_1195 , wr_751  , wr_447  );
  nor  g491( wr_1196 , wr_754  , wr_389  );
  nor  g492( wr_1217 , wr_751  , wr_778  );
  nor  g493( wr_1218 , wr_754  , wr_776  );
  nor  g494( wr_1451 , wr_743  , wr_447  );
  nor  g495( wr_1472 , wr_743  , wr_66   );
  nor  g496( wr_1300 , wr_743  , wr_847  );
  nor  g497( wr_1321 , wr_743  , wr_59   );
  nor  g498( wr_1380 , wr_743  , wr_27   );
  nor  g499( wr_1408 , wr_737  , wr_847  );
  nor  g500( wr_752  , wr_751  , wr_44   );
  nor  g501( wr_755  , wr_754  , wr_41   );
  nor  g502( wr_781  , wr_751  , wr_780  );
  nor  g503( wr_783  , wr_754  , wr_782  );
  nor  g504( wr_842  , wr_737  , wr_44   );
  nor  g505( wr_866  , wr_737  , wr_66   );
  nor  g506( wr_1044 , wr_748  , wr_389  );
  nor  g507( wr_1067 , wr_748  , wr_348  );
  nor  g508( wr_1126 , wr_751  , wr_389  );
  nor  g509( wr_1127 , wr_754  , wr_44   );
  nor  g510( wr_1149 , wr_751  , wr_782  );
  nor  g511( wr_1150 , wr_754  , wr_778  );
  nor  g512( wr_1194 , wr_748  , wr_44   );
  nor  g513( wr_1216 , wr_748  , wr_303  );
  nor  g514( wr_1450 , wr_737  , wr_389  );
  nor  g515( wr_1471 , wr_737  , wr_59   );
  nor  g516( wr_738  , wr_737  , wr_27   );
  nor  g517( wr_1123 , wr_737  , wr_47   );
  nor  g518( wr_1299 , wr_737  , wr_447  );
  nor  g519( wr_749  , wr_748  , wr_50   );
  nor  g520( wr_779  , wr_748  , wr_778  );
  nor  g521( wr_1043 , wr_743  , wr_44   );
  nor  g522( wr_1066 , wr_743  , wr_199  );
  nor  g523( wr_1125 , wr_748  , wr_41   );
  nor  g524( wr_1148 , wr_748  , wr_776  );
  nor  g525( wr_1193 , wr_743  , wr_41   );
  nor  g526( wr_1215 , wr_743  , wr_348  );
  nor  g527( wr_744  , wr_743  , wr_47   );
  nor  g528( wr_777  , wr_743  , wr_776  );
  nor  g529( wr_1042 , wr_737  , wr_41   );
  nor  g530( wr_1065 , wr_737  , wr_63   );
  nor  g531( wr_1124 , wr_743  , wr_50   );
  nor  g532( wr_1147 , wr_743  , wr_303  );
  nor  g533( wr_1192 , wr_737  , wr_50   );
  nor  g534( wr_1214 , wr_737  , wr_199  );
  nor  g535( wr_1404 , wr_726  , wr_389  );
  nor  g536( wr_775  , wr_737  , wr_303  );
  nor  g537( wr_838  , wr_726  , wr_50   );
  nor  g538( wr_864  , wr_726  , wr_27   );
  nor  g539( wr_1039 , wr_726  , wr_47   );
  nor  g540( wr_1146 , wr_737  , wr_348  );
  nor  g541( wr_1378 , wr_726  , wr_41   );
  not  g542( wr_1110 ,           wr_1109 );
  nor  g543( wr_1295 , wr_726  , wr_44   );
  not  g544( wr_699  ,           wr_698  );
  nor  g545( wr_727  , wr_726  , wr_66   );
  nor  g546( wr_1062 , wr_726  , wr_59   );
  nor  g547( wr_1105 , wr_110  , wr_184  );
  nor  g548( wr_704  , wr_703  , wr_702  );
  nor  g549( wr_837  , wr_836  , G77     );
  nor  g550( wr_1034 , wr_701  , wr_98   );
  nor  g551( wr_1185 , wr_701  , wr_124  );
  nor  g552( wr_1447 , wr_836  , G68     );
  nor  g553( wr_771  , wr_726  , wr_199  );
  nor  g554( wr_1143 , wr_726  , wr_63   );
  nor  g555( wr_1294 , wr_836  , G58     );
  nor  g556( wr_1375 , wr_836  , G50     );
  nor  g557( wr_696  , wr_695  , wr_29   );
  not  g558( wr_811  ,           wr_810  );
  nor  g559( wr_1103 , wr_695  , wr_669  );
  not  g560( wr_58   ,           wr_57   );
  not  g561( wr_74   ,           wr_73   );
  not  g562( wr_677  ,           wr_676  );
  nor  g563( wr_680  , wr_679  , wr_84   );
  nor  g564( wr_965  , wr_964  , wr_959  );
  nor  g565( wr_137  , wr_136  , wr_124  );
  nor  g566( wr_139  , wr_135  , wr_138  );
  nor  g567( wr_111  , wr_110  , wr_98   );
  nor  g568( wr_113  , wr_109  , wr_112  );
  nor  g569( wr_156  , wr_155  , wr_59   );
  nor  g570( wr_173  , wr_172  , wr_152  );
  nor  g571( wr_208  , wr_207  , wr_204  );
  nor  g572( wr_234  , wr_155  , wr_27   );
  nor  g573( wr_265  , wr_264  , wr_261  );
  nor  g574( wr_288  , wr_155  , wr_63   );
  nor  g575( wr_310  , wr_309  , wr_308  );
  nor  g576( wr_333  , wr_155  , wr_66   );
  nor  g577( wr_355  , wr_354  , wr_353  );
  nor  g578( wr_385  , wr_155  , wr_41   );
  nor  g579( wr_399  , wr_398  , wr_152  );
  nor  g580( wr_420  , wr_419  , wr_416  );
  nor  g581( wr_443  , wr_155  , wr_44   );
  nor  g582( wr_466  , wr_465  , wr_464  );
  nor  g583( wr_489  , wr_155  , wr_47   );
  nor  g584( wr_510  , wr_509  , wr_508  );
  nor  g585( wr_533  , wr_155  , wr_50   );
  nor  g586( wr_554  , wr_553  , wr_552  );
  nor  g587( wr_1413 , wr_1412 , wr_1411 );
  nor  g588( wr_849  , wr_848  , wr_846  );
  nor  g589( wr_871  , wr_870  , wr_869  );
  nor  g590( wr_1455 , wr_1454 , wr_1453 );
  nor  g591( wr_1476 , wr_1475 , wr_1474 );
  nor  g592( wr_1305 , wr_1304 , wr_1303 );
  nor  g593( wr_1325 , wr_1324 , wr_1323 );
  nor  g594( wr_1384 , wr_1383 , wr_1382 );
  nor  g595( wr_1047 , wr_1046 , wr_1045 );
  nor  g596( wr_1070 , wr_1069 , wr_1068 );
  nor  g597( wr_1197 , wr_1196 , wr_1195 );
  nor  g598( wr_1219 , wr_1218 , wr_1217 );
  nor  g599( wr_756  , wr_755  , wr_752  );
  nor  g600( wr_784  , wr_783  , wr_781  );
  nor  g601( wr_1128 , wr_1127 , wr_1126 );
  nor  g602( wr_1151 , wr_1150 , wr_1149 );
  nor  g603( wr_1111 , wr_1110 , wr_1106 );
  nor  g604( wr_1033 , wr_699  , G87     );
  nor  g605( wr_1184 , wr_699  , G97     );
  not  g606( wr_705  ,           wr_704  );
  nor  g607( wr_700  , wr_699  , G116    );
  nor  g608( wr_1104 , wr_699  , G107    );
  nor  g609( wr_75   , wr_74   , wr_58   );
  nor  g610( wr_678  , wr_677  , wr_670  );
  nor  g611( wr_140  , wr_139  , wr_137  );
  nor  g612( G358    , wr_113  , wr_111  );
  not  g613( wr_157  ,           wr_156  );
  not  g614( wr_209  ,           wr_208  );
  not  g615( wr_235  ,           wr_234  );
  not  g616( wr_266  ,           wr_265  );
  not  g617( wr_289  ,           wr_288  );
  not  g618( wr_311  ,           wr_310  );
  not  g619( wr_334  ,           wr_333  );
  not  g620( wr_356  ,           wr_355  );
  not  g621( wr_386  ,           wr_385  );
  not  g622( wr_421  ,           wr_420  );
  not  g623( wr_444  ,           wr_443  );
  not  g624( wr_467  ,           wr_466  );
  not  g625( wr_490  ,           wr_489  );
  not  g626( wr_511  ,           wr_510  );
  not  g627( wr_534  ,           wr_533  );
  not  g628( wr_555  ,           wr_554  );
  not  g629( wr_1414 ,           wr_1413 );
  not  g630( wr_850  ,           wr_849  );
  not  g631( wr_872  ,           wr_871  );
  not  g632( wr_1456 ,           wr_1455 );
  not  g633( wr_1477 ,           wr_1476 );
  not  g634( wr_1306 ,           wr_1305 );
  not  g635( wr_1326 ,           wr_1325 );
  not  g636( wr_1385 ,           wr_1384 );
  not  g637( wr_1048 ,           wr_1047 );
  not  g638( wr_1071 ,           wr_1070 );
  not  g639( wr_1198 ,           wr_1197 );
  not  g640( wr_1220 ,           wr_1219 );
  not  g641( wr_757  ,           wr_756  );
  not  g642( wr_785  ,           wr_784  );
  not  g643( wr_1129 ,           wr_1128 );
  not  g644( wr_1152 ,           wr_1151 );
  not  g645( wr_1112 ,           wr_1111 );
  nor  g646( wr_1035 , wr_1034 , wr_1033 );
  nor  g647( wr_1186 , wr_1185 , wr_1184 );
  nor  g648( wr_706  , wr_705  , wr_701  );
  nor  g649( wr_80   , wr_79   , wr_75   );
  nor  g650( wr_681  , wr_680  , wr_678  );
  not  g651( G351    ,           wr_140  );
  nor  g652( wr_158  , wr_157  , wr_147  );
  nor  g653( wr_210  , wr_209  , wr_191  );
  nor  g654( wr_236  , wr_235  , wr_147  );
  nor  g655( wr_267  , wr_266  , wr_254  );
  nor  g656( wr_290  , wr_289  , wr_147  );
  nor  g657( wr_312  , wr_311  , wr_191  );
  nor  g658( wr_335  , wr_334  , wr_147  );
  nor  g659( wr_357  , wr_356  , wr_191  );
  nor  g660( wr_387  , wr_386  , wr_384  );
  nor  g661( wr_422  , wr_421  , wr_408  );
  nor  g662( wr_445  , wr_444  , wr_384  );
  nor  g663( wr_468  , wr_467  , wr_408  );
  nor  g664( wr_491  , wr_490  , wr_384  );
  nor  g665( wr_512  , wr_511  , wr_408  );
  nor  g666( wr_535  , wr_534  , wr_384  );
  nor  g667( wr_556  , wr_555  , wr_408  );
  nor  g668( wr_1415 , wr_1414 , wr_1410 );
  nor  g669( wr_851  , wr_850  , wr_844  );
  nor  g670( wr_873  , wr_872  , wr_868  );
  nor  g671( wr_1457 , wr_1456 , wr_1452 );
  nor  g672( wr_1478 , wr_1477 , wr_1473 );
  nor  g673( wr_1307 , wr_1306 , wr_1301 );
  nor  g674( wr_1327 , wr_1326 , wr_1322 );
  nor  g675( wr_1386 , wr_1385 , wr_1381 );
  nor  g676( wr_1049 , wr_1048 , wr_1044 );
  nor  g677( wr_1072 , wr_1071 , wr_1067 );
  nor  g678( wr_1199 , wr_1198 , wr_1194 );
  nor  g679( wr_1221 , wr_1220 , wr_1216 );
  nor  g680( wr_758  , wr_757  , wr_749  );
  nor  g681( wr_786  , wr_785  , wr_779  );
  nor  g682( wr_1130 , wr_1129 , wr_1125 );
  nor  g683( wr_1153 , wr_1152 , wr_1148 );
  nor  g684( wr_1113 , wr_1112 , G45     );
  not  g685( wr_1036 ,           wr_1035 );
  not  g686( wr_1187 ,           wr_1186 );
  nor  g687( wr_707  , wr_706  , wr_700  );
  nor  g688( wr_86   , wr_85   , wr_80   );
  not  g689( wr_682  ,           wr_681  );
  nor  g690( wr_174  , wr_173  , wr_158  );
  nor  g691( wr_211  , wr_210  , wr_177  );
  not  g692( wr_215  ,           wr_210  );
  nor  g693( wr_223  , wr_210  , wr_222  );
  nor  g694( wr_247  , wr_246  , wr_236  );
  nor  g695( wr_268  , wr_267  , wr_177  );
  not  g696( wr_271  ,           wr_267  );
  nor  g697( wr_278  , wr_267  , wr_222  );
  nor  g698( wr_298  , wr_297  , wr_290  );
  nor  g699( wr_313  , wr_312  , wr_177  );
  not  g700( wr_316  ,           wr_312  );
  nor  g701( wr_323  , wr_312  , wr_222  );
  nor  g702( wr_343  , wr_342  , wr_335  );
  nor  g703( wr_358  , wr_357  , wr_177  );
  not  g704( wr_361  ,           wr_357  );
  nor  g705( wr_368  , wr_357  , wr_222  );
  nor  g706( wr_400  , wr_399  , wr_387  );
  nor  g707( wr_423  , wr_422  , wr_177  );
  not  g708( wr_426  ,           wr_422  );
  nor  g709( wr_433  , wr_422  , wr_222  );
  nor  g710( wr_454  , wr_453  , wr_445  );
  nor  g711( wr_469  , wr_468  , wr_177  );
  not  g712( wr_472  ,           wr_468  );
  nor  g713( wr_479  , wr_468  , wr_222  );
  nor  g714( wr_499  , wr_498  , wr_491  );
  nor  g715( wr_513  , wr_512  , wr_177  );
  not  g716( wr_516  ,           wr_512  );
  nor  g717( wr_523  , wr_512  , wr_222  );
  nor  g718( wr_543  , wr_542  , wr_535  );
  nor  g719( wr_557  , wr_556  , wr_177  );
  not  g720( wr_560  ,           wr_556  );
  nor  g721( wr_567  , wr_556  , wr_222  );
  nor  g722( wr_647  , wr_312  , G179    );
  not  g723( wr_1416 ,           wr_1415 );
  not  g724( wr_852  ,           wr_851  );
  not  g725( wr_874  ,           wr_873  );
  not  g726( wr_1458 ,           wr_1457 );
  not  g727( wr_1479 ,           wr_1478 );
  not  g728( wr_1308 ,           wr_1307 );
  not  g729( wr_1328 ,           wr_1327 );
  not  g730( wr_1387 ,           wr_1386 );
  not  g731( wr_1050 ,           wr_1049 );
  not  g732( wr_1073 ,           wr_1072 );
  not  g733( wr_1200 ,           wr_1199 );
  not  g734( wr_1222 ,           wr_1221 );
  not  g735( wr_759  ,           wr_758  );
  not  g736( wr_787  ,           wr_786  );
  not  g737( wr_1131 ,           wr_1130 );
  not  g738( wr_1154 ,           wr_1153 );
  nor  g739( wr_1114 , wr_1113 , wr_1105 );
  nor  g740( wr_1037 , wr_1036 , wr_694  );
  nor  g741( wr_1188 , wr_1187 , wr_694  );
  not  g742( wr_708  ,           wr_707  );
  not  g743( wr_87   ,           wr_86   );
  not  g744( wr_175  ,           wr_174  );
  not  g745( wr_212  ,           wr_211  );
  nor  g746( wr_216  , wr_215  , wr_214  );
  not  g747( wr_224  ,           wr_223  );
  nor  g748( wr_227  , wr_215  , wr_226  );
  not  g749( wr_248  ,           wr_247  );
  not  g750( wr_269  ,           wr_268  );
  nor  g751( wr_272  , wr_271  , wr_214  );
  not  g752( wr_279  ,           wr_278  );
  nor  g753( wr_281  , wr_271  , wr_226  );
  not  g754( wr_299  ,           wr_298  );
  not  g755( wr_314  ,           wr_313  );
  nor  g756( wr_317  , wr_316  , wr_214  );
  not  g757( wr_324  ,           wr_323  );
  nor  g758( wr_326  , wr_316  , wr_226  );
  not  g759( wr_344  ,           wr_343  );
  not  g760( wr_359  ,           wr_358  );
  nor  g761( wr_362  , wr_361  , wr_214  );
  not  g762( wr_369  ,           wr_368  );
  nor  g763( wr_371  , wr_361  , wr_226  );
  not  g764( wr_401  ,           wr_400  );
  not  g765( wr_424  ,           wr_423  );
  nor  g766( wr_427  , wr_426  , wr_214  );
  not  g767( wr_434  ,           wr_433  );
  nor  g768( wr_436  , wr_426  , wr_226  );
  not  g769( wr_455  ,           wr_454  );
  not  g770( wr_470  ,           wr_469  );
  nor  g771( wr_473  , wr_472  , wr_214  );
  not  g772( wr_480  ,           wr_479  );
  nor  g773( wr_482  , wr_472  , wr_226  );
  not  g774( wr_500  ,           wr_499  );
  not  g775( wr_514  ,           wr_513  );
  nor  g776( wr_517  , wr_516  , wr_214  );
  not  g777( wr_524  ,           wr_523  );
  nor  g778( wr_526  , wr_516  , wr_226  );
  not  g779( wr_544  ,           wr_543  );
  not  g780( wr_558  ,           wr_557  );
  nor  g781( wr_561  , wr_560  , wr_214  );
  not  g782( wr_568  ,           wr_567  );
  nor  g783( wr_570  , wr_560  , wr_226  );
  not  g784( wr_648  ,           wr_647  );
  nor  g785( wr_1417 , wr_1416 , wr_1409 );
  nor  g786( wr_853  , wr_852  , wr_843  );
  nor  g787( wr_875  , wr_874  , wr_867  );
  nor  g788( wr_1459 , wr_1458 , wr_1451 );
  nor  g789( wr_1480 , wr_1479 , wr_1472 );
  nor  g790( wr_1309 , wr_1308 , wr_1300 );
  nor  g791( wr_1329 , wr_1328 , wr_1321 );
  nor  g792( wr_1388 , wr_1387 , wr_1380 );
  nor  g793( wr_1051 , wr_1050 , wr_1043 );
  nor  g794( wr_1074 , wr_1073 , wr_1066 );
  nor  g795( wr_1201 , wr_1200 , wr_1193 );
  nor  g796( wr_1223 , wr_1222 , wr_1215 );
  nor  g797( wr_760  , wr_759  , wr_744  );
  nor  g798( wr_788  , wr_787  , wr_777  );
  nor  g799( wr_1132 , wr_1131 , wr_1124 );
  nor  g800( wr_1155 , wr_1154 , wr_1147 );
  not  g801( wr_1115 ,           wr_1114 );
  nor  g802( wr_1038 , wr_1037 , wr_715  );
  nor  g803( wr_1189 , wr_1188 , wr_715  );
  nor  g804( wr_709  , wr_708  , wr_696  );
  nor  g805( G361    , wr_87   , wr_40   );
  nor  g806( wr_176  , wr_175  , wr_145  );
  not  g807( wr_217  ,           wr_216  );
  nor  g808( wr_249  , wr_248  , wr_233  );
  not  g809( wr_273  ,           wr_272  );
  nor  g810( wr_300  , wr_299  , wr_287  );
  not  g811( wr_318  ,           wr_317  );
  nor  g812( wr_345  , wr_344  , wr_332  );
  not  g813( wr_363  ,           wr_362  );
  nor  g814( wr_402  , wr_401  , wr_383  );
  not  g815( wr_428  ,           wr_427  );
  nor  g816( wr_456  , wr_455  , wr_442  );
  not  g817( wr_474  ,           wr_473  );
  nor  g818( wr_501  , wr_500  , wr_488  );
  not  g819( wr_518  ,           wr_517  );
  nor  g820( wr_545  , wr_544  , wr_532  );
  not  g821( wr_562  ,           wr_561  );
  nor  g822( wr_649  , wr_648  , wr_357  );
  not  g823( wr_1418 ,           wr_1417 );
  not  g824( wr_854  ,           wr_853  );
  not  g825( wr_876  ,           wr_875  );
  not  g826( wr_1460 ,           wr_1459 );
  not  g827( wr_1481 ,           wr_1480 );
  not  g828( wr_1310 ,           wr_1309 );
  not  g829( wr_1330 ,           wr_1329 );
  not  g830( wr_1389 ,           wr_1388 );
  not  g831( wr_1052 ,           wr_1051 );
  not  g832( wr_1075 ,           wr_1074 );
  not  g833( wr_1202 ,           wr_1201 );
  not  g834( wr_1224 ,           wr_1223 );
  not  g835( wr_761  ,           wr_760  );
  not  g836( wr_789  ,           wr_788  );
  not  g837( wr_1133 ,           wr_1132 );
  not  g838( wr_1156 ,           wr_1155 );
  nor  g839( wr_1116 , wr_1115 , wr_701  );
  nor  g840( wr_716  , wr_715  , wr_709  );
  nor  g841( wr_213  , wr_212  , wr_176  );
  nor  g842( wr_218  , wr_217  , wr_176  );
  not  g843( wr_221  ,           wr_176  );
  nor  g844( wr_270  , wr_269  , wr_249  );
  nor  g845( wr_274  , wr_273  , wr_249  );
  not  g846( wr_277  ,           wr_249  );
  nor  g847( wr_315  , wr_314  , wr_300  );
  nor  g848( wr_319  , wr_318  , wr_300  );
  not  g849( wr_322  ,           wr_300  );
  nor  g850( wr_360  , wr_359  , wr_345  );
  nor  g851( wr_364  , wr_363  , wr_345  );
  not  g852( wr_367  ,           wr_345  );
  nor  g853( wr_425  , wr_424  , wr_402  );
  nor  g854( wr_429  , wr_428  , wr_402  );
  not  g855( wr_432  ,           wr_402  );
  nor  g856( wr_471  , wr_470  , wr_456  );
  nor  g857( wr_475  , wr_474  , wr_456  );
  not  g858( wr_478  ,           wr_456  );
  nor  g859( wr_515  , wr_514  , wr_501  );
  nor  g860( wr_519  , wr_518  , wr_501  );
  not  g861( wr_522  ,           wr_501  );
  nor  g862( wr_559  , wr_558  , wr_545  );
  nor  g863( wr_563  , wr_562  , wr_545  );
  not  g864( wr_566  ,           wr_545  );
  nor  g865( wr_819  , wr_623  , wr_501  );
  nor  g866( wr_902  , wr_901  , wr_402  );
  nor  g867( wr_654  , wr_361  , wr_318  );
  nor  g868( wr_907  , wr_623  , wr_545  );
  not  g869( wr_650  ,           wr_649  );
  nor  g870( wr_969  , wr_623  , wr_176  );
  nor  g871( wr_1419 , wr_1418 , wr_1408 );
  nor  g872( wr_855  , wr_854  , wr_842  );
  nor  g873( wr_877  , wr_876  , wr_866  );
  nor  g874( wr_1461 , wr_1460 , wr_1450 );
  nor  g875( wr_1482 , wr_1481 , wr_1471 );
  nor  g876( wr_624  , wr_623  , wr_345  );
  nor  g877( wr_1311 , wr_1310 , wr_1299 );
  nor  g878( wr_1331 , wr_1330 , wr_738  );
  nor  g879( wr_1390 , wr_1389 , wr_1123 );
  nor  g880( wr_1353 , wr_901  , wr_456  );
  nor  g881( wr_634  , wr_623  , wr_300  );
  nor  g882( wr_1053 , wr_1052 , wr_1042 );
  nor  g883( wr_1076 , wr_1075 , wr_1065 );
  nor  g884( wr_1203 , wr_1202 , wr_1192 );
  nor  g885( wr_1225 , wr_1224 , wr_1214 );
  nor  g886( wr_980  , wr_623  , wr_249  );
  nor  g887( wr_762  , wr_761  , wr_738  );
  nor  g888( wr_790  , wr_789  , wr_775  );
  nor  g889( wr_1134 , wr_1133 , wr_1123 );
  nor  g890( wr_1157 , wr_1156 , wr_1146 );
  nor  g891( wr_1117 , wr_1116 , wr_1104 );
  nor  g892( wr_219  , wr_218  , wr_213  );
  nor  g893( wr_225  , wr_224  , wr_221  );
  nor  g894( wr_228  , wr_227  , wr_221  );
  nor  g895( wr_275  , wr_274  , wr_270  );
  nor  g896( wr_280  , wr_279  , wr_277  );
  nor  g897( wr_282  , wr_281  , wr_277  );
  nor  g898( wr_320  , wr_319  , wr_315  );
  nor  g899( wr_327  , wr_326  , wr_322  );
  nor  g900( wr_365  , wr_364  , wr_360  );
  nor  g901( wr_370  , wr_369  , wr_367  );
  nor  g902( wr_372  , wr_371  , wr_367  );
  nor  g903( wr_437  , wr_436  , wr_432  );
  nor  g904( wr_476  , wr_475  , wr_471  );
  nor  g905( wr_481  , wr_480  , wr_478  );
  nor  g906( wr_483  , wr_482  , wr_478  );
  nor  g907( wr_520  , wr_519  , wr_515  );
  nor  g908( wr_525  , wr_524  , wr_522  );
  nor  g909( wr_527  , wr_526  , wr_522  );
  nor  g910( wr_564  , wr_563  , wr_559  );
  nor  g911( wr_569  , wr_568  , wr_566  );
  nor  g912( wr_571  , wr_570  , wr_566  );
  nor  g913( wr_325  , wr_324  , wr_322  );
  nor  g914( wr_430  , wr_429  , wr_425  );
  nor  g915( wr_435  , wr_434  , wr_432  );
  not  g916( wr_820  ,           wr_819  );
  not  g917( wr_903  ,           wr_902  );
  not  g918( wr_655  ,           wr_654  );
  not  g919( wr_908  ,           wr_907  );
  nor  g920( wr_651  , wr_650  , wr_267  );
  not  g921( wr_970  ,           wr_969  );
  not  g922( wr_1420 ,           wr_1419 );
  not  g923( wr_856  ,           wr_855  );
  not  g924( wr_878  ,           wr_877  );
  not  g925( wr_1462 ,           wr_1461 );
  not  g926( wr_1483 ,           wr_1482 );
  not  g927( wr_625  ,           wr_624  );
  not  g928( wr_1312 ,           wr_1311 );
  not  g929( wr_1332 ,           wr_1331 );
  not  g930( wr_1391 ,           wr_1390 );
  not  g931( wr_1354 ,           wr_1353 );
  not  g932( wr_635  ,           wr_634  );
  not  g933( wr_1054 ,           wr_1053 );
  not  g934( wr_1077 ,           wr_1076 );
  not  g935( wr_1204 ,           wr_1203 );
  not  g936( wr_1226 ,           wr_1225 );
  not  g937( wr_981  ,           wr_980  );
  not  g938( wr_763  ,           wr_762  );
  not  g939( wr_791  ,           wr_790  );
  not  g940( wr_1135 ,           wr_1134 );
  not  g941( wr_1158 ,           wr_1157 );
  not  g942( wr_1118 ,           wr_1117 );
  not  g943( wr_220  ,           wr_219  );
  not  g944( wr_229  ,           wr_228  );
  not  g945( wr_276  ,           wr_275  );
  not  g946( wr_283  ,           wr_282  );
  not  g947( wr_366  ,           wr_365  );
  not  g948( wr_373  ,           wr_372  );
  not  g949( wr_477  ,           wr_476  );
  not  g950( wr_484  ,           wr_483  );
  not  g951( wr_521  ,           wr_520  );
  not  g952( wr_528  ,           wr_527  );
  not  g953( wr_565  ,           wr_564  );
  not  g954( wr_572  ,           wr_571  );
  not  g955( wr_328  ,           wr_327  );
  not  g956( wr_438  ,           wr_437  );
  not  g957( wr_321  ,           wr_320  );
  not  g958( wr_431  ,           wr_430  );
  nor  g959( wr_936  , wr_621  , wr_520  );
  nor  g960( wr_656  , wr_655  , wr_271  );
  not  g961( wr_652  ,           wr_651  );
  nor  g962( wr_629  , wr_621  , wr_320  );
  nor  g963( wr_1421 , wr_1420 , wr_1407 );
  nor  g964( wr_857  , wr_856  , wr_841  );
  nor  g965( wr_879  , wr_878  , wr_735  );
  nor  g966( wr_927  , wr_621  , wr_564  );
  nor  g967( wr_930  , wr_900  , wr_430  );
  nor  g968( wr_1463 , wr_1462 , wr_1449 );
  nor  g969( wr_1484 , wr_1483 , wr_1122 );
  nor  g970( wr_1313 , wr_1312 , wr_1298 );
  nor  g971( wr_1333 , wr_1332 , wr_1191 );
  nor  g972( wr_1392 , wr_1391 , wr_1041 );
  nor  g973( wr_622  , wr_621  , wr_365  );
  nor  g974( wr_990  , wr_621  , wr_219  );
  nor  g975( wr_1055 , wr_1054 , wr_1041 );
  nor  g976( wr_1078 , wr_1077 , wr_1064 );
  nor  g977( wr_1205 , wr_1204 , wr_1191 );
  nor  g978( wr_1227 , wr_1226 , wr_1213 );
  nor  g979( wr_764  , wr_763  , wr_735  );
  nor  g980( wr_792  , wr_791  , wr_774  );
  nor  g981( wr_1136 , wr_1135 , wr_1122 );
  nor  g982( wr_1159 , wr_1158 , wr_1145 );
  nor  g983( wr_1119 , wr_1118 , wr_1103 );
  nor  g984( wr_230  , wr_229  , wr_225  );
  nor  g985( wr_284  , wr_283  , wr_280  );
  nor  g986( wr_374  , wr_373  , wr_370  );
  nor  g987( wr_485  , wr_484  , wr_481  );
  nor  g988( wr_529  , wr_528  , wr_525  );
  nor  g989( wr_573  , wr_572  , wr_569  );
  nor  g990( wr_329  , wr_328  , wr_325  );
  nor  g991( wr_439  , wr_438  , wr_435  );
  not  g992( wr_937  ,           wr_936  );
  not  g993( wr_657  ,           wr_656  );
  nor  g994( wr_653  , wr_652  , wr_210  );
  not  g995( wr_630  ,           wr_629  );
  not  g996( wr_1422 ,           wr_1421 );
  not  g997( wr_858  ,           wr_857  );
  not  g998( wr_880  ,           wr_879  );
  not  g999( wr_928  ,           wr_927  );
  not g1000( wr_1464 ,           wr_1463 );
  not g1001( wr_1485 ,           wr_1484 );
  not g1002( wr_1314 ,           wr_1313 );
  not g1003( wr_1334 ,           wr_1333 );
  not g1004( wr_1393 ,           wr_1392 );
  not g1005( wr_985  ,           wr_622  );
  not g1006( wr_1056 ,           wr_1055 );
  not g1007( wr_1079 ,           wr_1078 );
  not g1008( wr_1206 ,           wr_1205 );
  not g1009( wr_1228 ,           wr_1227 );
  not g1010( wr_765  ,           wr_764  );
  not g1011( wr_793  ,           wr_792  );
  not g1012( wr_1137 ,           wr_1136 );
  not g1013( wr_1160 ,           wr_1159 );
  nor g1014( wr_1120 , wr_1119 , wr_715  );
  nor g1015( wr_231  , wr_230  , wr_220  );
  nor g1016( wr_285  , wr_284  , wr_276  );
  nor g1017( wr_375  , wr_374  , wr_366  );
  nor g1018( wr_486  , wr_485  , wr_477  );
  nor g1019( wr_530  , wr_529  , wr_521  );
  nor g1020( wr_574  , wr_573  , wr_565  );
  nor g1021( wr_330  , wr_329  , wr_321  );
  nor g1022( wr_440  , wr_439  , wr_431  );
  nor g1023( wr_658  , wr_657  , wr_215  );
  nor g1024( wr_1423 , wr_1422 , wr_1406 );
  nor g1025( wr_859  , wr_858  , wr_840  );
  nor g1026( wr_881  , wr_880  , wr_865  );
  nor g1027( wr_1465 , wr_1464 , wr_1448 );
  nor g1028( wr_1486 , wr_1485 , wr_1470 );
  nor g1029( wr_1315 , wr_1314 , wr_1297 );
  nor g1030( wr_1335 , wr_1334 , wr_1320 );
  nor g1031( wr_1394 , wr_1393 , wr_1379 );
  nor g1032( wr_1057 , wr_1056 , wr_1040 );
  nor g1033( wr_1080 , wr_1079 , wr_1063 );
  nor g1034( wr_1207 , wr_1206 , wr_1190 );
  nor g1035( wr_1229 , wr_1228 , wr_1212 );
  nor g1036( wr_766  , wr_765  , wr_732  );
  nor g1037( wr_794  , wr_793  , wr_773  );
  nor g1038( wr_1138 , wr_1137 , wr_1121 );
  nor g1039( wr_1161 , wr_1160 , wr_1144 );
  not g1040( wr_232  ,           wr_231  );
  not g1041( wr_286  ,           wr_285  );
  not g1042( wr_376  ,           wr_375  );
  not g1043( wr_487  ,           wr_486  );
  not g1044( wr_531  ,           wr_530  );
  not g1045( wr_575  ,           wr_574  );
  nor g1046( wr_821  , wr_820  , wr_530  );
  not g1047( wr_331  ,           wr_330  );
  not g1048( wr_441  ,           wr_440  );
  nor g1049( wr_904  , wr_903  , wr_440  );
  nor g1050( wr_909  , wr_908  , wr_574  );
  nor g1051( wr_659  , wr_658  , wr_653  );
  nor g1052( wr_971  , wr_970  , wr_231  );
  nor g1053( wr_626  , wr_625  , wr_375  );
  nor g1054( wr_1355 , wr_1354 , wr_486  );
  not g1055( wr_1424 ,           wr_1423 );
  nor g1056( wr_636  , wr_635  , wr_330  );
  not g1057( wr_860  ,           wr_859  );
  not g1058( wr_882  ,           wr_881  );
  not g1059( wr_1466 ,           wr_1465 );
  not g1060( wr_1487 ,           wr_1486 );
  not g1061( wr_1316 ,           wr_1315 );
  not g1062( wr_1336 ,           wr_1335 );
  not g1063( wr_1395 ,           wr_1394 );
  nor g1064( wr_982  , wr_981  , wr_285  );
  not g1065( wr_1058 ,           wr_1057 );
  not g1066( wr_1081 ,           wr_1080 );
  not g1067( wr_1208 ,           wr_1207 );
  not g1068( wr_1230 ,           wr_1229 );
  not g1069( wr_767  ,           wr_766  );
  not g1070( wr_795  ,           wr_794  );
  not g1071( wr_1139 ,           wr_1138 );
  not g1072( wr_1162 ,           wr_1161 );
  nor g1073( wr_583  , wr_376  , wr_286  );
  nor g1074( wr_588  , wr_365  , wr_286  );
  nor g1075( wr_582  , wr_286  , wr_219  );
  nor g1076( wr_598  , wr_575  , wr_487  );
  nor g1077( wr_822  , wr_819  , wr_531  );
  nor g1078( wr_377  , wr_376  , wr_331  );
  nor g1079( wr_603  , wr_564  , wr_487  );
  nor g1080( wr_905  , wr_902  , wr_441  );
  nor g1081( wr_576  , wr_575  , wr_531  );
  nor g1082( wr_910  , wr_907  , wr_575  );
  nor g1083( wr_972  , wr_969  , wr_232  );
  nor g1084( wr_597  , wr_487  , wr_430  );
  nor g1085( wr_660  , wr_659  , wr_623  );
  nor g1086( wr_627  , wr_624  , wr_376  );
  nor g1087( wr_1356 , wr_1353 , wr_487  );
  nor g1088( wr_637  , wr_634  , wr_331  );
  nor g1089( wr_1425 , wr_1424 , wr_1404 );
  nor g1090( wr_861  , wr_860  , wr_838  );
  nor g1091( wr_883  , wr_882  , wr_864  );
  nor g1092( wr_1467 , wr_1466 , wr_1378 );
  nor g1093( wr_1488 , wr_1487 , wr_1039 );
  nor g1094( wr_983  , wr_980  , wr_286  );
  nor g1095( wr_1317 , wr_1316 , wr_1295 );
  nor g1096( wr_1337 , wr_1336 , wr_838  );
  nor g1097( wr_1396 , wr_1395 , wr_1378 );
  nor g1098( wr_1059 , wr_1058 , wr_1039 );
  nor g1099( wr_1082 , wr_1081 , wr_1062 );
  nor g1100( wr_1209 , wr_1208 , wr_864  );
  nor g1101( wr_1231 , wr_1230 , wr_727  );
  nor g1102( wr_768  , wr_767  , wr_727  );
  nor g1103( wr_796  , wr_795  , wr_771  );
  nor g1104( wr_1140 , wr_1139 , wr_1062 );
  nor g1105( wr_1163 , wr_1162 , wr_1143 );
  not g1106( wr_584  ,           wr_583  );
  not g1107( wr_589  ,           wr_588  );
  not g1108( wr_599  ,           wr_598  );
  nor g1109( wr_823  , wr_822  , wr_821  );
  not g1110( wr_378  ,           wr_377  );
  not g1111( wr_604  ,           wr_603  );
  nor g1112( wr_906  , wr_905  , wr_904  );
  not g1113( wr_577  ,           wr_576  );
  nor g1114( wr_911  , wr_910  , wr_909  );
  nor g1115( wr_973  , wr_972  , wr_971  );
  nor g1116( wr_628  , wr_627  , wr_626  );
  nor g1117( wr_1357 , wr_1356 , wr_1355 );
  nor g1118( wr_638  , wr_637  , wr_636  );
  not g1119( wr_1426 ,           wr_1425 );
  not g1120( wr_862  ,           wr_861  );
  not g1121( wr_884  ,           wr_883  );
  not g1122( wr_1468 ,           wr_1467 );
  not g1123( wr_1489 ,           wr_1488 );
  nor g1124( wr_984  , wr_983  , wr_982  );
  not g1125( wr_1318 ,           wr_1317 );
  not g1126( wr_1338 ,           wr_1337 );
  not g1127( wr_1397 ,           wr_1396 );
  not g1128( wr_1060 ,           wr_1059 );
  not g1129( wr_1083 ,           wr_1082 );
  not g1130( wr_1210 ,           wr_1209 );
  not g1131( wr_1232 ,           wr_1231 );
  not g1132( wr_769  ,           wr_768  );
  not g1133( wr_797  ,           wr_796  );
  not g1134( wr_1141 ,           wr_1140 );
  not g1135( wr_1164 ,           wr_1163 );
  nor g1136( wr_585  , wr_584  , wr_320  );
  nor g1137( wr_590  , wr_589  , wr_232  );
  nor g1138( wr_600  , wr_599  , wr_520  );
  nor g1139( wr_379  , wr_378  , wr_286  );
  nor g1140( wr_605  , wr_604  , wr_441  );
  nor g1141( wr_938  , wr_937  , wr_906  );
  nor g1142( wr_578  , wr_577  , wr_487  );
  nor g1143( wr_912  , wr_911  , wr_823  );
  nor g1144( wr_987  , wr_973  , wr_630  );
  nor g1145( wr_929  , wr_928  , wr_906  );
  not g1146( wr_1359 ,           wr_1357 );
  nor g1147( wr_974  , wr_973  , wr_638  );
  nor g1148( wr_986  , wr_973  , wr_985  );
  nor g1149( wr_1251 , wr_937  , wr_911  );
  not g1150( wr_1275 ,           wr_911  );
  nor g1151( wr_1427 , wr_1426 , wr_1403 );
  nor g1152( wr_863  , wr_862  , G33     );
  nor g1153( wr_885  , wr_884  , wr_146  );
  nor g1154( wr_1469 , wr_1468 , G33     );
  nor g1155( wr_1490 , wr_1489 , wr_146  );
  not g1156( wr_826  ,           wr_823  );
  not g1157( wr_996  ,           wr_984  );
  not g1158( wr_1260 ,           wr_906  );
  nor g1159( wr_1319 , wr_1318 , G33     );
  nor g1160( wr_1339 , wr_1338 , wr_146  );
  nor g1161( wr_1398 , wr_1397 , wr_1377 );
  nor g1162( wr_631  , wr_630  , wr_628  );
  not g1163( wr_1017 ,           wr_628  );
  nor g1164( wr_639  , wr_638  , wr_628  );
  not g1165( wr_1007 ,           wr_973  );
  nor g1166( wr_1016 , wr_629  , wr_628  );
  nor g1167( wr_1061 , wr_1060 , G33     );
  nor g1168( wr_1084 , wr_1083 , wr_146  );
  nor g1169( wr_1211 , wr_1210 , G33     );
  nor g1170( wr_1233 , wr_1232 , wr_146  );
  nor g1171( wr_1014 , wr_638  , wr_641  );
  nor g1172( wr_770  , wr_769  , G33     );
  nor g1173( wr_798  , wr_797  , wr_146  );
  nor g1174( wr_1142 , wr_1141 , G33     );
  nor g1175( wr_1165 , wr_1164 , wr_146  );
  not g1176( wr_685  ,           wr_638  );
  nor g1177( wr_684  , wr_638  , G330    );
  not g1178( wr_586  ,           wr_585  );
  not g1179( wr_601  ,           wr_600  );
  not g1180( wr_380  ,           wr_379  );
  not g1181( wr_939  ,           wr_938  );
  not g1182( wr_579  ,           wr_578  );
  not g1183( wr_913  ,           wr_912  );
  not g1184( wr_988  ,           wr_987  );
  not g1185( wr_975  ,           wr_974  );
  nor g1186( wr_1428 , wr_1427 , wr_1402 );
  nor g1187( wr_886  , wr_885  , wr_863  );
  nor g1188( wr_1491 , wr_1490 , wr_1469 );
  nor g1189( wr_1340 , wr_1339 , wr_1319 );
  nor g1190( wr_632  , wr_631  , wr_622  );
  nor g1191( wr_834  , wr_826  , wr_690  );
  nor g1192( wr_1018 , wr_630  , wr_1017 );
  nor g1193( wr_1446 , wr_1275 , wr_690  );
  not g1194( wr_640  ,           wr_639  );
  nor g1195( wr_1085 , wr_1084 , wr_1061 );
  nor g1196( wr_1234 , wr_1233 , wr_1211 );
  nor g1197( wr_1293 , wr_1260 , wr_690  );
  nor g1198( wr_1374 , wr_1359 , wr_690  );
  not g1199( wr_1015 ,           wr_1014 );
  nor g1200( wr_799  , wr_798  , wr_770  );
  nor g1201( wr_1166 , wr_1165 , wr_1142 );
  nor g1202( wr_1032 , wr_996  , wr_692  );
  nor g1203( wr_1183 , wr_1007 , wr_692  );
  nor g1204( wr_693  , wr_692  , wr_685  );
  nor g1205( wr_1102 , wr_692  , wr_1017 );
  nor g1206( wr_686  , wr_685  , wr_641  );
  nor g1207( wr_587  , wr_586  , wr_232  );
  nor g1208( wr_602  , wr_601  , wr_441  );
  nor g1209( wr_381  , wr_380  , wr_232  );
  nor g1210( wr_940  , wr_939  , wr_911  );
  nor g1211( wr_580  , wr_579  , wr_441  );
  nor g1212( wr_989  , wr_988  , wr_628  );
  nor g1213( wr_976  , wr_975  , wr_628  );
  not g1214( wr_1429 ,           wr_1428 );
  nor g1215( wr_887  , wr_886  , wr_717  );
  nor g1216( wr_1492 , wr_1491 , wr_717  );
  nor g1217( wr_1341 , wr_1340 , wr_717  );
  not g1218( wr_633  ,           wr_632  );
  nor g1219( wr_1008 , wr_1007 , wr_632  );
  nor g1220( wr_1019 , wr_1018 , wr_1016 );
  nor g1221( wr_1004 , wr_640  , wr_641  );
  nor g1222( wr_1086 , wr_1085 , wr_717  );
  nor g1223( wr_1235 , wr_1234 , wr_717  );
  nor g1224( wr_800  , wr_799  , wr_717  );
  nor g1225( wr_1167 , wr_1166 , wr_717  );
  nor g1226( wr_687  , wr_686  , wr_684  );
  nor g1227( wr_591  , wr_590  , wr_587  );
  nor g1228( wr_606  , wr_605  , wr_602  );
  not g1229( wr_382  ,           wr_381  );
  not g1230( wr_581  ,           wr_580  );
  nor g1231( wr_991  , wr_990  , wr_989  );
  not g1232( wr_977  ,           wr_976  );
  nor g1233( wr_1430 , wr_1429 , wr_1398 );
  nor g1234( wr_888  , wr_887  , wr_837  );
  nor g1235( wr_1493 , wr_1492 , wr_1447 );
  nor g1236( wr_1342 , wr_1341 , wr_1294 );
  nor g1237( wr_1006 , wr_973  , wr_633  );
  not g1238( wr_1020 ,           wr_1019 );
  not g1239( wr_1005 ,           wr_1004 );
  nor g1240( wr_1022 , wr_1019 , wr_1014 );
  nor g1241( wr_1087 , wr_1086 , wr_1038 );
  nor g1242( wr_1236 , wr_1235 , wr_1189 );
  nor g1243( wr_801  , wr_800  , wr_716  );
  nor g1244( wr_1168 , wr_1167 , wr_1120 );
  nor g1245( wr_813  , wr_808  , wr_687  );
  nor g1246( wr_688  , wr_687  , wr_679  );
  nor g1247( wr_642  , wr_633  , wr_641  );
  not g1248( wr_592  ,           wr_591  );
  not g1249( wr_607  ,           wr_606  );
  nor g1250( wr_661  , wr_621  , wr_382  );
  not g1251( wr_992  ,           wr_991  );
  nor g1252( wr_978  , wr_977  , wr_641  );
  nor g1253( wr_1431 , wr_1430 , wr_717  );
  not g1254( wr_889  ,           wr_888  );
  not g1255( wr_1494 ,           wr_1493 );
  not g1256( wr_1343 ,           wr_1342 );
  nor g1257( wr_1009 , wr_1008 , wr_1006 );
  nor g1258( wr_1021 , wr_1020 , wr_1015 );
  not g1259( wr_1088 ,           wr_1087 );
  not g1260( wr_1237 ,           wr_1236 );
  not g1261( wr_802  ,           wr_801  );
  not g1262( wr_1169 ,           wr_1168 );
  not g1263( wr_643  ,           wr_642  );
  nor g1264( G372    , wr_581  , wr_382  );
  nor g1265( wr_593  , wr_592  , wr_276  );
  nor g1266( wr_608  , wr_607  , wr_477  );
  nor g1267( wr_662  , wr_661  , wr_660  );
  nor g1268( wr_993  , wr_992  , wr_986  );
  not g1269( wr_979  ,           wr_978  );
  nor g1270( wr_1432 , wr_1431 , wr_1375 );
  nor g1271( wr_890  , wr_889  , wr_834  );
  nor g1272( wr_1495 , wr_1494 , wr_1446 );
  nor g1273( wr_1344 , wr_1343 , wr_1293 );
  not g1274( wr_1010 ,           wr_1009 );
  nor g1275( wr_1012 , wr_1009 , wr_1004 );
  nor g1276( wr_1023 , wr_1022 , wr_1021 );
  nor g1277( wr_1089 , wr_1088 , wr_1032 );
  nor g1278( wr_1238 , wr_1237 , wr_1183 );
  nor g1279( wr_803  , wr_802  , wr_693  );
  nor g1280( wr_1170 , wr_1169 , wr_1102 );
  nor g1281( wr_644  , wr_643  , wr_640  );
  not g1282( wr_594  ,           wr_593  );
  not g1283( wr_609  ,           wr_608  );
  nor g1284( wr_914  , wr_913  , wr_662  );
  nor g1285( wr_918  , wr_662  , wr_581  );
  nor g1286( wr_1245 , wr_911  , wr_662  );
  nor g1287( wr_1268 , wr_823  , wr_662  );
  not g1288( wr_994  ,           wr_993  );
  nor g1289( wr_997  , wr_993  , wr_996  );
  nor g1290( wr_817  , wr_662  , wr_641  );
  not g1291( wr_1433 ,           wr_1432 );
  not g1292( wr_891  ,           wr_890  );
  not g1293( wr_1496 ,           wr_1495 );
  not g1294( wr_1345 ,           wr_1344 );
  nor g1295( wr_1011 , wr_1010 , wr_1005 );
  not g1296( wr_1090 ,           wr_1089 );
  not g1297( wr_1239 ,           wr_1238 );
  not g1298( wr_1097 ,           wr_1023 );
  not g1299( wr_804  ,           wr_803  );
  not g1300( wr_1171 ,           wr_1170 );
  nor g1301( wr_1173 , wr_1023 , wr_808  );
  nor g1302( wr_645  , wr_644  , wr_633  );
  nor g1303( wr_595  , wr_594  , wr_582  );
  nor g1304( wr_610  , wr_609  , wr_597  );
  not g1305( wr_915  ,           wr_914  );
  not g1306( wr_920  ,           wr_918  );
  not g1307( wr_1246 ,           wr_1245 );
  not g1308( wr_1269 ,           wr_1268 );
  nor g1309( wr_995  , wr_994  , wr_984  );
  not g1310( wr_818  ,           wr_817  );
  nor g1311( wr_1434 , wr_1433 , wr_1374 );
  nor g1312( wr_892  , wr_891  , wr_811  );
  nor g1313( wr_1497 , wr_1496 , wr_811  );
  nor g1314( wr_1346 , wr_1345 , wr_811  );
  nor g1315( wr_1013 , wr_1012 , wr_1011 );
  nor g1316( wr_1091 , wr_1090 , wr_811  );
  nor g1317( wr_1240 , wr_1239 , wr_811  );
  nor g1318( wr_812  , wr_811  , wr_804  );
  nor g1319( wr_1172 , wr_1171 , wr_811  );
  not g1320( G399    ,           wr_645  );
  nor g1321( wr_646  , wr_621  , wr_595  );
  not g1322( wr_611  ,           wr_610  );
  nor g1323( wr_916  , wr_915  , wr_906  );
  nor g1324( wr_1247 , wr_1246 , wr_823  );
  nor g1325( wr_1270 , wr_1269 , wr_641  );
  nor g1326( wr_998  , wr_997  , wr_995  );
  not g1327( wr_1435 ,           wr_1434 );
  not g1328( wr_1177 ,           wr_1013 );
  nor g1329( wr_1241 , wr_1013 , wr_808  );
  nor g1330( wr_814  , wr_813  , wr_812  );
  nor g1331( wr_1174 , wr_1173 , wr_1172 );
  nor g1332( wr_596  , wr_595  , wr_581  );
  not g1333( wr_825  ,           wr_646  );
  not g1334( wr_917  ,           wr_916  );
  nor g1335( wr_663  , wr_646  , wr_641  );
  nor g1336( wr_824  , wr_823  , wr_646  );
  not g1337( wr_1248 ,           wr_1247 );
  not g1338( wr_1271 ,           wr_1270 );
  not g1339( wr_999  ,           wr_998  );
  nor g1340( wr_1001 , wr_998  , wr_978  );
  nor g1341( wr_1436 , wr_1435 , wr_811  );
  nor g1342( wr_1242 , wr_1241 , wr_1240 );
  not g1343( wr_815  ,           wr_814  );
  not g1344( wr_1175 ,           wr_1174 );
  nor g1345( wr_921  , wr_920  , wr_916  );
  nor g1346( wr_612  , wr_611  , wr_596  );
  nor g1347( wr_931  , wr_823  , wr_825  );
  nor g1348( wr_1252 , wr_911  , wr_825  );
  nor g1349( wr_925  , wr_825  , wr_581  );
  nor g1350( wr_1351 , wr_917  , wr_641  );
  nor g1351( wr_827  , wr_826  , wr_825  );
  not g1352( wr_664  ,           wr_663  );
  nor g1353( wr_1249 , wr_1248 , wr_641  );
  nor g1354( wr_1000 , wr_999  , wr_979  );
  not g1355( wr_1243 ,           wr_1242 );
  nor g1356( wr_816  , wr_815  , wr_688  );
  nor g1357( wr_919  , wr_918  , wr_917  );
  not g1358( G369    ,           wr_612  );
  not g1359( wr_932  ,           wr_931  );
  not g1360( wr_1253 ,           wr_1252 );
  nor g1361( wr_926  , wr_925  , wr_611  );
  nor g1362( wr_1272 , wr_936  , wr_931  );
  not g1363( wr_1352 ,           wr_1351 );
  nor g1364( wr_828  , wr_827  , wr_824  );
  nor g1365( wr_665  , wr_664  , wr_662  );
  not g1366( wr_1250 ,           wr_1249 );
  nor g1367( wr_1002 , wr_1001 , wr_1000 );
  not g1368( G396    ,           wr_816  );
  nor g1369( wr_922  , wr_921  , wr_919  );
  nor g1370( wr_933  , wr_932  , wr_906  );
  nor g1371( wr_1254 , wr_1253 , wr_823  );
  not g1372( wr_948  ,           wr_926  );
  not g1373( wr_1273 ,           wr_1272 );
  nor g1374( wr_1276 , wr_1272 , wr_1275 );
  not g1375( wr_829  ,           wr_828  );
  nor g1376( wr_666  , wr_665  , wr_646  );
  nor g1377( wr_831  , wr_828  , wr_817  );
  nor g1378( wr_1092 , wr_1002 , wr_808  );
  nor g1379( wr_923  , wr_922  , wr_641  );
  not g1380( wr_934  ,           wr_933  );
  nor g1381( wr_1255 , wr_1254 , wr_927  );
  nor g1382( wr_1282 , wr_948  , wr_641  );
  nor g1383( wr_1274 , wr_1273 , wr_911  );
  nor g1384( wr_830  , wr_829  , wr_818  );
  not g1385( wr_1024 ,           wr_666  );
  nor g1386( wr_1003 , wr_1002 , wr_666  );
  nor g1387( wr_1093 , wr_1092 , wr_1091 );
  nor g1388( wr_1098 , wr_1097 , wr_666  );
  not g1389( wr_924  ,           wr_923  );
  nor g1390( wr_667  , wr_666  , G1      );
  nor g1391( wr_935  , wr_934  , wr_911  );
  not g1392( wr_1256 ,           wr_1255 );
  not g1393( wr_1283 ,           wr_1282 );
  nor g1394( wr_1277 , wr_1276 , wr_1274 );
  nor g1395( wr_832  , wr_831  , wr_830  );
  nor g1396( wr_1025 , wr_1002 , wr_1024 );
  nor g1397( wr_1096 , wr_1023 , wr_1024 );
  not g1398( wr_1094 ,           wr_1093 );
  nor g1399( wr_683  , wr_682  , wr_667  );
  nor g1400( wr_941  , wr_940  , wr_935  );
  nor g1401( wr_1257 , wr_1256 , wr_1251 );
  nor g1402( wr_1284 , wr_1283 , wr_920  );
  not g1403( wr_1278 ,           wr_1277 );
  nor g1404( wr_1280 , wr_1277 , wr_1270 );
  nor g1405( wr_893  , wr_832  , wr_808  );
  not g1406( wr_1026 ,           wr_1025 );
  nor g1407( wr_833  , wr_832  , wr_679  );
  not g1408( wr_1178 ,           wr_1096 );
  nor g1409( wr_1180 , wr_1096 , wr_1013 );
  nor g1410( wr_1099 , wr_1098 , wr_1096 );
  not g1411( G364    ,           wr_683  );
  not g1412( wr_942  ,           wr_941  );
  not g1413( wr_1258 ,           wr_1257 );
  nor g1414( wr_1261 , wr_1257 , wr_1260 );
  nor g1415( wr_1285 , wr_1284 , wr_948  );
  nor g1416( wr_1279 , wr_1278 , wr_1271 );
  nor g1417( wr_894  , wr_893  , wr_892  );
  nor g1418( wr_1027 , wr_1026 , wr_1023 );
  nor g1419( wr_1179 , wr_1178 , wr_1177 );
  not g1420( wr_1100 ,           wr_1099 );
  nor g1421( wr_943  , wr_942  , wr_930  );
  nor g1422( wr_1259 , wr_1258 , wr_906  );
  not g1423( wr_1286 ,           wr_1285 );
  nor g1424( wr_1281 , wr_1280 , wr_1279 );
  not g1425( wr_895  ,           wr_894  );
  not g1426( wr_1028 ,           wr_1027 );
  nor g1427( wr_1181 , wr_1180 , wr_1179 );
  nor g1428( wr_1101 , wr_1100 , wr_679  );
  not g1429( wr_944  ,           wr_943  );
  nor g1430( wr_1262 , wr_1261 , wr_1259 );
  not g1431( wr_1441 ,           wr_1281 );
  nor g1432( wr_1287 , wr_1286 , wr_1281 );
  nor g1433( wr_1498 , wr_1281 , wr_808  );
  nor g1434( wr_896  , wr_895  , wr_833  );
  nor g1435( wr_1029 , wr_1028 , wr_1013 );
  nor g1436( wr_1182 , wr_1181 , wr_679  );
  nor g1437( wr_1176 , wr_1175 , wr_1101 );
  nor g1438( wr_945  , wr_944  , wr_929  );
  not g1439( wr_1263 ,           wr_1262 );
  nor g1440( wr_1265 , wr_1262 , wr_1249 );
  nor g1441( wr_1442 , wr_1285 , wr_1441 );
  not g1442( wr_1288 ,           wr_1287 );
  nor g1443( wr_1499 , wr_1498 , wr_1497 );
  not g1444( G384    ,           wr_896  );
  nor g1445( wr_1030 , wr_1029 , wr_1003 );
  nor g1446( wr_1244 , wr_1243 , wr_1182 );
  not g1447( G393    ,           wr_1176 );
  nor g1448( wr_1526 , wr_1176 , G396    );
  not g1449( wr_946  ,           wr_945  );
  nor g1450( wr_1360 , wr_1359 , wr_945  );
  nor g1451( wr_1264 , wr_1263 , wr_1250 );
  nor g1452( wr_1443 , wr_1442 , wr_1287 );
  not g1453( wr_1500 ,           wr_1499 );
  nor g1454( wr_1031 , wr_1030 , wr_679  );
  not g1455( G390    ,           wr_1244 );
  nor g1456( wr_949  , wr_945  , wr_948  );
  nor g1457( wr_1527 , G393    , wr_816  );
  nor g1458( wr_1358 , wr_1357 , wr_946  );
  nor g1459( wr_1266 , wr_1265 , wr_1264 );
  not g1460( wr_1444 ,           wr_1443 );
  nor g1461( wr_1095 , wr_1094 , wr_1031 );
  nor g1462( wr_947  , wr_946  , wr_926  );
  nor g1463( wr_1528 , wr_1527 , wr_1526 );
  nor g1464( wr_1361 , wr_1360 , wr_1358 );
  not g1465( wr_1267 ,           wr_1266 );
  nor g1466( wr_1290 , wr_1287 , wr_1266 );
  nor g1467( wr_1347 , wr_1266 , wr_808  );
  nor g1468( wr_1445 , wr_1444 , wr_679  );
  not g1469( G387    ,           wr_1095 );
  nor g1470( wr_950  , wr_949  , wr_947  );
  nor g1471( wr_1523 , G390    , wr_1095 );
  not g1472( wr_1529 ,           wr_1528 );
  not g1473( wr_1362 ,           wr_1361 );
  nor g1474( wr_1364 , wr_1361 , wr_1351 );
  nor g1475( wr_1289 , wr_1288 , wr_1267 );
  nor g1476( wr_1348 , wr_1347 , wr_1346 );
  nor g1477( wr_1501 , wr_1500 , wr_1445 );
  nor g1478( wr_1502 , G390    , G387    );
  nor g1479( wr_1524 , wr_1244 , G387    );
  not g1480( wr_951  ,           wr_950  );
  nor g1481( wr_953  , wr_950  , wr_923  );
  nor g1482( wr_1363 , wr_1362 , wr_1352 );
  nor g1483( wr_1291 , wr_1290 , wr_1289 );
  not g1484( wr_1349 ,           wr_1348 );
  not g1485( G381    ,           wr_1501 );
  nor g1486( wr_1545 , wr_1501 , G384    );
  not g1487( wr_1503 ,           wr_1502 );
  nor g1488( wr_1525 , wr_1524 , wr_1523 );
  nor g1489( wr_952  , wr_951  , wr_924  );
  nor g1490( wr_1365 , wr_1364 , wr_1363 );
  nor g1491( wr_1292 , wr_1291 , wr_679  );
  nor g1492( wr_1546 , G381    , wr_896  );
  nor g1493( wr_1504 , wr_1503 , G396    );
  not g1494( wr_1531 ,           wr_1525 );
  nor g1495( wr_954  , wr_953  , wr_952  );
  nor g1496( wr_1530 , wr_1529 , wr_1525 );
  nor g1497( wr_1367 , wr_1365 , wr_1286 );
  nor g1498( wr_1366 , wr_1365 , wr_1285 );
  nor g1499( wr_1437 , wr_1365 , wr_808  );
  nor g1500( wr_1350 , wr_1349 , wr_1292 );
  nor g1501( wr_1547 , wr_1546 , wr_1545 );
  not g1502( wr_1505 ,           wr_1504 );
  nor g1503( wr_1532 , wr_1528 , wr_1531 );
  nor g1504( wr_958  , wr_957  , wr_954  );
  not g1505( wr_1368 ,           wr_1367 );
  nor g1506( wr_1438 , wr_1437 , wr_1436 );
  nor g1507( wr_1535 , wr_1515 , wr_1350 );
  not g1508( wr_1555 ,           wr_1547 );
  not g1509( G378    ,           wr_1350 );
  nor g1510( wr_1552 , wr_1547 , wr_1551 );
  nor g1511( wr_1548 , wr_1547 , wr_1544 );
  nor g1512( wr_1506 , wr_1505 , G393    );
  nor g1513( wr_1533 , wr_1532 , wr_1530 );
  nor g1514( wr_966  , wr_965  , wr_958  );
  nor g1515( wr_1369 , wr_1368 , wr_1281 );
  not g1516( wr_1439 ,           wr_1438 );
  not g1517( wr_1536 ,           wr_1535 );
  nor g1518( wr_1556 , wr_1555 , wr_1551 );
  nor g1519( wr_1559 , wr_1555 , wr_1544 );
  not g1520( wr_1553 ,           wr_1552 );
  nor g1521( wr_1517 , wr_1516 , G378    );
  not g1522( wr_1549 ,           wr_1548 );
  not g1523( wr_1507 ,           wr_1506 );
  not g1524( wr_1534 ,           wr_1533 );
  not g1525( wr_967  ,           wr_966  );
  not g1526( wr_1370 ,           wr_1369 );
  not g1527( wr_1557 ,           wr_1556 );
  not g1528( wr_1560 ,           wr_1559 );
  not g1529( wr_1518 ,           wr_1517 );
  nor g1530( wr_968  , wr_967  , wr_899  );
  nor g1531( wr_1371 , wr_1370 , wr_1266 );
  not g1532( G367    ,           wr_968  );
  nor g1533( wr_1372 , wr_1371 , wr_1366 );
  nor g1534( wr_1373 , wr_1372 , wr_679  );
  nor g1535( wr_1440 , wr_1439 , wr_1373 );
  nor g1536( wr_1537 , wr_1515 , wr_1440 );
  not g1537( G375    ,           wr_1440 );
  nor g1538( wr_1571 , wr_1440 , G378    );
  not g1539( wr_1539 ,           wr_1537 );
  nor g1540( wr_1538 , wr_1537 , wr_1536 );
  nor g1541( wr_1508 , G375    , G378    );
  nor g1542( wr_1572 , G375    , wr_1350 );
  nor g1543( wr_1519 , wr_1518 , G375    );
  nor g1544( wr_1540 , wr_1539 , wr_1535 );
  not g1545( wr_1509 ,           wr_1508 );
  nor g1546( wr_1573 , wr_1572 , wr_1571 );
  nor g1547( wr_1541 , wr_1540 , wr_1538 );
  nor g1548( wr_1510 , wr_1509 , G384    );
  not g1549( wr_1575 ,           wr_1573 );
  nor g1550( wr_1574 , wr_1573 , wr_1555 );
  not g1551( wr_1542 ,           wr_1541 );
  nor g1552( wr_1561 , wr_1560 , wr_1541 );
  not g1553( wr_1511 ,           wr_1510 );
  nor g1554( wr_1554 , wr_1553 , wr_1541 );
  nor g1555( wr_1576 , wr_1575 , wr_1547 );
  nor g1556( wr_1558 , wr_1557 , wr_1542 );
  nor g1557( wr_1512 , wr_1511 , G381    );
  nor g1558( wr_1550 , wr_1549 , wr_1542 );
  nor g1559( wr_1577 , wr_1576 , wr_1574 );
  nor g1560( wr_1562 , wr_1561 , wr_1558 );
  not g1561( wr_1513 ,           wr_1512 );
  not g1562( wr_1579 ,           wr_1577 );
  nor g1563( wr_1578 , wr_1577 , wr_1534 );
  not g1564( wr_1563 ,           wr_1562 );
  nor g1565( wr_1514 , wr_1513 , wr_1507 );
  nor g1566( wr_1580 , wr_1579 , wr_1533 );
  nor g1567( wr_1564 , wr_1563 , wr_1554 );
  nor g1568( wr_1520 , wr_1519 , wr_1514 );
  not g1569( G407    ,           wr_1514 );
  nor g1570( G402    , wr_1580 , wr_1578 );
  not g1571( wr_1565 ,           wr_1564 );
  not g1572( wr_1521 ,           wr_1520 );
  nor g1573( wr_1566 , wr_1565 , wr_1550 );
  nor g1574( wr_1522 , wr_1521 , wr_613  );
  not g1575( wr_1567 ,           wr_1566 );
  nor g1576( wr_1569 , wr_1566 , wr_1533 );
  not g1577( G409    ,           wr_1522 );
  nor g1578( wr_1568 , wr_1567 , wr_1534 );
  nor g1579( wr_1570 , wr_1569 , wr_1568 );
  not g1580( G405    ,           wr_1570 );

endmodule
