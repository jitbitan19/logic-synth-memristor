// NOR_NOT mapped module b07_C

module b07_C (
  input  STATO_REG_0__SCAN_IN,
  input  STATO_REG_1__SCAN_IN,
  input  PUNTI_RETTA_REG_7__SCAN_IN,
  input  PUNTI_RETTA_REG_6__SCAN_IN,
  input  PUNTI_RETTA_REG_5__SCAN_IN,
  input  PUNTI_RETTA_REG_4__SCAN_IN,
  input  PUNTI_RETTA_REG_3__SCAN_IN,
  input  PUNTI_RETTA_REG_2__SCAN_IN,
  input  PUNTI_RETTA_REG_1__SCAN_IN,
  input  PUNTI_RETTA_REG_0__SCAN_IN,
  input  CONT_REG_7__SCAN_IN,
  input  CONT_REG_6__SCAN_IN,
  input  CONT_REG_5__SCAN_IN,
  input  CONT_REG_4__SCAN_IN,
  input  CONT_REG_3__SCAN_IN,
  input  CONT_REG_2__SCAN_IN,
  input  CONT_REG_1__SCAN_IN,
  input  CONT_REG_0__SCAN_IN,
  input  MAR_REG_7__SCAN_IN,
  input  MAR_REG_6__SCAN_IN,
  input  MAR_REG_5__SCAN_IN,
  input  MAR_REG_4__SCAN_IN,
  input  MAR_REG_3__SCAN_IN,
  input  MAR_REG_2__SCAN_IN,
  input  MAR_REG_1__SCAN_IN,
  input  MAR_REG_0__SCAN_IN,
  input  X_REG_7__SCAN_IN,
  input  X_REG_6__SCAN_IN,
  input  X_REG_5__SCAN_IN,
  input  X_REG_4__SCAN_IN,
  input  X_REG_3__SCAN_IN,
  input  X_REG_2__SCAN_IN,
  input  X_REG_1__SCAN_IN,
  input  X_REG_0__SCAN_IN,
  input  Y_REG_3__SCAN_IN,
  input  Y_REG_1__SCAN_IN,
  input  Y_REG_5__SCAN_IN,
  input  T_REG_3__SCAN_IN,
  input  T_REG_5__SCAN_IN,
  input  T_REG_1__SCAN_IN,
  input  T_REG_0__SCAN_IN,
  input  T_REG_4__SCAN_IN,
  input  T_REG_6__SCAN_IN,
  input  T_REG_2__SCAN_IN,
  input  Y_REG_4__SCAN_IN,
  input  Y_REG_0__SCAN_IN,
  input  Y_REG_2__SCAN_IN,
  input  Y_REG_6__SCAN_IN,
  input  STATO_REG_2__SCAN_IN,
  output PUNTI_RETTA_7_,
  output PUNTI_RETTA_6_,
  output PUNTI_RETTA_5_,
  output PUNTI_RETTA_4_,
  output PUNTI_RETTA_3_,
  output PUNTI_RETTA_2_,
  output PUNTI_RETTA_1_,
  output PUNTI_RETTA_0_,
  output PUNTI_RETTA_REG_7__SCAN_OUT,
  output PUNTI_RETTA_REG_6__SCAN_OUT,
  output PUNTI_RETTA_REG_5__SCAN_OUT,
  output PUNTI_RETTA_REG_4__SCAN_OUT,
  output PUNTI_RETTA_REG_3__SCAN_OUT,
  output PUNTI_RETTA_REG_2__SCAN_OUT,
  output PUNTI_RETTA_REG_1__SCAN_OUT,
  output PUNTI_RETTA_REG_0__SCAN_OUT,
  output CONT_REG_7__SCAN_OUT,
  output CONT_REG_6__SCAN_OUT,
  output CONT_REG_5__SCAN_OUT,
  output CONT_REG_4__SCAN_OUT,
  output CONT_REG_3__SCAN_OUT,
  output CONT_REG_2__SCAN_OUT,
  output CONT_REG_1__SCAN_OUT,
  output CONT_REG_0__SCAN_OUT,
  output MAR_REG_7__SCAN_OUT,
  output MAR_REG_6__SCAN_OUT,
  output MAR_REG_5__SCAN_OUT,
  output MAR_REG_4__SCAN_OUT,
  output MAR_REG_3__SCAN_OUT,
  output MAR_REG_2__SCAN_OUT,
  output MAR_REG_1__SCAN_OUT,
  output MAR_REG_0__SCAN_OUT,
  output X_REG_7__SCAN_OUT,
  output X_REG_6__SCAN_OUT,
  output X_REG_5__SCAN_OUT,
  output X_REG_4__SCAN_OUT,
  output X_REG_3__SCAN_OUT,
  output X_REG_2__SCAN_OUT,
  output X_REG_1__SCAN_OUT,
  output X_REG_0__SCAN_OUT,
  output Y_REG_3__SCAN_OUT,
  output Y_REG_1__SCAN_OUT,
  output Y_REG_5__SCAN_OUT,
  output T_REG_3__SCAN_OUT,
  output T_REG_5__SCAN_OUT,
  output T_REG_1__SCAN_OUT,
  output T_REG_0__SCAN_OUT,
  output T_REG_4__SCAN_OUT,
  output T_REG_6__SCAN_OUT,
  output T_REG_2__SCAN_OUT,
  output Y_REG_4__SCAN_OUT,
  output Y_REG_0__SCAN_OUT,
  output Y_REG_2__SCAN_OUT,
  output Y_REG_6__SCAN_OUT,
  output STATO_REG_2__SCAN_OUT,
  output STATO_REG_1__SCAN_OUT,
  output STATO_REG_0__SCAN_OUT);

  wire wr_58;
  wire wr_59;
  wire wr_60;
  wire wr_61;
  wire wr_62;
  wire wr_63;
  wire wr_64;
  wire wr_65;
  wire wr_66;
  wire wr_67;
  wire wr_68;
  wire wr_69;
  wire wr_70;
  wire wr_71;
  wire wr_72;
  wire wr_73;
  wire wr_74;
  wire wr_75;
  wire wr_76;
  wire wr_77;
  wire wr_78;
  wire wr_79;
  wire wr_80;
  wire wr_81;
  wire wr_82;
  wire wr_83;
  wire wr_84;
  wire wr_85;
  wire wr_86;
  wire wr_87;
  wire wr_88;
  wire wr_89;
  wire wr_90;
  wire wr_91;
  wire wr_92;
  wire wr_93;
  wire wr_94;
  wire wr_95;
  wire wr_96;
  wire wr_97;
  wire wr_98;
  wire wr_99;
  wire wr_100;
  wire wr_101;
  wire wr_102;
  wire wr_103;
  wire wr_104;
  wire wr_105;
  wire wr_106;
  wire wr_107;
  wire wr_108;
  wire wr_109;
  wire wr_110;
  wire wr_111;
  wire wr_112;
  wire wr_113;
  wire wr_114;
  wire wr_115;
  wire wr_116;
  wire wr_117;
  wire wr_118;
  wire wr_119;
  wire wr_120;
  wire wr_121;
  wire wr_122;
  wire wr_123;
  wire wr_124;
  wire wr_125;
  wire wr_126;
  wire wr_127;
  wire wr_128;
  wire wr_129;
  wire wr_130;
  wire wr_131;
  wire wr_132;
  wire wr_133;
  wire wr_134;
  wire wr_135;
  wire wr_136;
  wire wr_137;
  wire wr_138;
  wire wr_139;
  wire wr_140;
  wire wr_141;
  wire wr_142;
  wire wr_143;
  wire wr_144;
  wire wr_145;
  wire wr_146;
  wire wr_147;
  wire wr_148;
  wire wr_149;
  wire wr_150;
  wire wr_151;
  wire wr_152;
  wire wr_153;
  wire wr_154;
  wire wr_155;
  wire wr_156;
  wire wr_157;
  wire wr_158;
  wire wr_159;
  wire wr_160;
  wire wr_161;
  wire wr_162;
  wire wr_163;
  wire wr_164;
  wire wr_165;
  wire wr_166;
  wire wr_167;
  wire wr_168;
  wire wr_169;
  wire wr_170;
  wire wr_171;
  wire wr_172;
  wire wr_173;
  wire wr_174;
  wire wr_175;
  wire wr_176;
  wire wr_177;
  wire wr_178;
  wire wr_179;
  wire wr_180;
  wire wr_181;
  wire wr_182;
  wire wr_183;
  wire wr_184;
  wire wr_185;
  wire wr_186;
  wire wr_187;
  wire wr_188;
  wire wr_189;
  wire wr_190;
  wire wr_191;
  wire wr_192;
  wire wr_193;
  wire wr_194;
  wire wr_195;
  wire wr_196;
  wire wr_197;
  wire wr_198;
  wire wr_199;
  wire wr_200;
  wire wr_201;
  wire wr_202;
  wire wr_203;
  wire wr_204;
  wire wr_205;
  wire wr_206;
  wire wr_207;
  wire wr_208;
  wire wr_209;
  wire wr_210;
  wire wr_211;
  wire wr_212;
  wire wr_213;
  wire wr_214;
  wire wr_215;
  wire wr_216;
  wire wr_217;
  wire wr_218;
  wire wr_219;
  wire wr_220;
  wire wr_221;
  wire wr_222;
  wire wr_223;
  wire wr_224;
  wire wr_225;
  wire wr_226;
  wire wr_227;
  wire wr_228;
  wire wr_229;
  wire wr_230;
  wire wr_231;
  wire wr_232;
  wire wr_233;
  wire wr_234;
  wire wr_235;
  wire wr_236;
  wire wr_237;
  wire wr_238;
  wire wr_239;
  wire wr_240;
  wire wr_241;
  wire wr_242;
  wire wr_243;
  wire wr_244;
  wire wr_245;
  wire wr_246;
  wire wr_247;
  wire wr_248;
  wire wr_249;
  wire wr_250;
  wire wr_251;
  wire wr_252;
  wire wr_253;
  wire wr_254;
  wire wr_255;
  wire wr_256;
  wire wr_257;
  wire wr_258;
  wire wr_259;
  wire wr_260;
  wire wr_261;
  wire wr_262;
  wire wr_263;
  wire wr_264;
  wire wr_265;
  wire wr_266;
  wire wr_267;
  wire wr_268;
  wire wr_269;
  wire wr_270;
  wire wr_271;
  wire wr_272;
  wire wr_273;
  wire wr_274;
  wire wr_275;
  wire wr_276;
  wire wr_277;
  wire wr_278;
  wire wr_279;
  wire wr_280;
  wire wr_281;
  wire wr_282;
  wire wr_283;
  wire wr_284;
  wire wr_285;
  wire wr_286;
  wire wr_287;
  wire wr_288;
  wire wr_289;
  wire wr_290;
  wire wr_291;
  wire wr_292;
  wire wr_293;
  wire wr_294;
  wire wr_295;
  wire wr_296;
  wire wr_297;
  wire wr_298;
  wire wr_299;
  wire wr_300;
  wire wr_301;
  wire wr_302;
  wire wr_303;
  wire wr_304;
  wire wr_305;
  wire wr_306;
  wire wr_307;
  wire wr_308;
  wire wr_309;
  wire wr_310;
  wire wr_311;
  wire wr_312;
  wire wr_313;
  wire wr_314;
  wire wr_315;
  wire wr_316;
  wire wr_317;
  wire wr_318;
  wire wr_319;
  wire wr_320;
  wire wr_321;
  wire wr_322;
  wire wr_323;
  wire wr_324;
  wire wr_325;
  wire wr_326;
  wire wr_327;
  wire wr_328;
  wire wr_329;
  wire wr_330;
  wire wr_331;
  wire wr_332;
  wire wr_333;
  wire wr_334;
  wire wr_335;
  wire wr_336;
  wire wr_337;
  wire wr_338;
  wire wr_339;
  wire wr_340;
  wire wr_341;
  wire wr_342;
  wire wr_343;
  wire wr_344;
  wire wr_345;
  wire wr_346;
  wire wr_347;
  wire wr_348;
  wire wr_349;
  wire wr_350;
  wire wr_351;
  wire wr_352;
  wire wr_353;
  wire wr_354;
  wire wr_355;
  wire wr_356;
  wire wr_357;
  wire wr_358;
  wire wr_359;
  wire wr_360;
  wire wr_361;
  wire wr_362;
  wire wr_363;
  wire wr_364;
  wire wr_365;
  wire wr_366;
  wire wr_367;
  wire wr_368;
  wire wr_369;
  wire wr_370;
  wire wr_371;
  wire wr_372;
  wire wr_373;
  wire wr_374;
  wire wr_375;
  wire wr_376;
  wire wr_377;
  wire wr_378;
  wire wr_379;
  wire wr_380;
  wire wr_381;
  wire wr_382;
  wire wr_383;
  wire wr_384;
  wire wr_385;
  wire wr_386;
  wire wr_387;
  wire wr_388;
  wire wr_389;
  wire wr_390;
  wire wr_391;
  wire wr_392;
  wire wr_393;
  wire wr_394;
  wire wr_395;
  wire wr_396;
  wire wr_397;
  wire wr_398;
  wire wr_399;
  wire wr_400;
  wire wr_401;
  wire wr_402;
  wire wr_403;
  wire wr_404;
  wire wr_405;
  wire wr_406;
  wire wr_407;
  wire wr_408;
  wire wr_409;
  wire wr_410;
  wire wr_411;
  wire wr_412;
  wire wr_413;
  wire wr_414;
  wire wr_415;
  wire wr_416;
  wire wr_417;
  wire wr_418;
  wire wr_419;
  wire wr_420;
  wire wr_421;
  wire wr_422;
  wire wr_423;
  wire wr_424;
  wire wr_425;
  wire wr_426;
  wire wr_427;
  wire wr_428;
  wire wr_429;
  wire wr_430;
  wire wr_431;
  wire wr_432;
  wire wr_433;
  wire wr_434;
  wire wr_435;
  wire wr_436;
  wire wr_437;
  wire wr_438;
  wire wr_439;
  wire wr_440;
  wire wr_441;
  wire wr_442;
  wire wr_443;
  wire wr_444;
  wire wr_445;
  wire wr_446;
  wire wr_447;
  wire wr_448;
  wire wr_449;
  wire wr_450;
  wire wr_451;
  wire wr_452;
  wire wr_453;
  wire wr_454;
  wire wr_455;
  wire wr_456;
  wire wr_457;
  wire wr_458;
  wire wr_459;
  wire wr_460;
  wire wr_461;
  wire wr_462;
  wire wr_463;
  wire wr_464;
  wire wr_465;
  wire wr_466;
  wire wr_467;
  wire wr_468;
  wire wr_469;
  wire wr_470;
  wire wr_471;
  wire wr_472;
  wire wr_473;
  wire wr_474;
  wire wr_475;
  wire wr_476;
  wire wr_477;
  wire wr_478;
  wire wr_479;
  wire wr_480;
  wire wr_481;
  wire wr_482;
  wire wr_483;
  wire wr_484;
  wire wr_485;
  wire wr_486;
  wire wr_487;
  wire wr_488;
  wire wr_489;
  wire wr_490;
  wire wr_491;
  wire wr_492;
  wire wr_493;
  wire wr_494;
  wire wr_495;
  wire wr_496;
  wire wr_497;
  wire wr_498;
  wire wr_499;
  wire wr_500;
  wire wr_501;
  wire wr_502;
  wire wr_503;
  wire wr_504;
  wire wr_505;
  wire wr_506;
  wire wr_507;
  wire wr_508;
  wire wr_509;
  wire wr_510;
  wire wr_511;
  wire wr_512;
  wire wr_513;
  wire wr_514;
  wire wr_515;
  wire wr_516;
  wire wr_517;
  wire wr_518;
  wire wr_519;
  wire wr_520;
  wire wr_521;
  wire wr_522;
  wire wr_523;
  wire wr_524;
  wire wr_525;
  wire wr_526;
  wire wr_527;
  wire wr_528;
  wire wr_529;
  wire wr_530;
  wire wr_531;
  wire wr_532;
  wire wr_533;
  wire wr_534;
  wire wr_535;
  wire wr_536;
  wire wr_537;
  wire wr_538;
  wire wr_539;
  wire wr_540;
  wire wr_541;
  wire wr_542;
  wire wr_543;
  wire wr_544;
  wire wr_545;
  wire wr_546;
  wire wr_547;
  wire wr_548;
  wire wr_549;
  wire wr_550;
  wire wr_551;
  wire wr_552;
  wire wr_553;
  wire wr_554;
  wire wr_555;
  wire wr_556;
  wire wr_557;
  wire wr_558;
  wire wr_559;
  wire wr_560;
  wire wr_561;

  not    g1( wr_59   ,           STATO_REG_1__SCAN_IN);
  not    g2( wr_60   ,           STATO_REG_2__SCAN_IN);
  not    g3( wr_82   ,           STATO_REG_0__SCAN_IN);
  nor    g4( wr_91   , STATO_REG_1__SCAN_IN, STATO_REG_0__SCAN_IN);
  not    g5( wr_122  ,           Y_REG_4__SCAN_IN);
  not    g6( wr_124  ,           T_REG_4__SCAN_IN);
  not    g7( wr_137  ,           X_REG_3__SCAN_IN);
  not    g8( wr_139  ,           Y_REG_3__SCAN_IN);
  not    g9( wr_141  ,           T_REG_3__SCAN_IN);
  not   g10( wr_147  ,           CONT_REG_3__SCAN_IN);
  not   g11( wr_154  ,           X_REG_2__SCAN_IN);
  not   g12( wr_156  ,           Y_REG_2__SCAN_IN);
  not   g13( wr_158  ,           T_REG_2__SCAN_IN);
  not   g14( wr_164  ,           CONT_REG_2__SCAN_IN);
  not   g15( wr_171  ,           X_REG_1__SCAN_IN);
  not   g16( wr_173  ,           Y_REG_1__SCAN_IN);
  not   g17( wr_175  ,           T_REG_1__SCAN_IN);
  not   g18( wr_181  ,           CONT_REG_1__SCAN_IN);
  not   g19( wr_185  ,           Y_REG_0__SCAN_IN);
  not   g20( wr_187  ,           X_REG_0__SCAN_IN);
  not   g21( wr_189  ,           T_REG_0__SCAN_IN);
  not   g22( wr_197  ,           CONT_REG_0__SCAN_IN);
  not   g23( wr_63   ,           MAR_REG_3__SCAN_IN);
  not   g24( wr_103  ,           Y_REG_5__SCAN_IN);
  not   g25( wr_106  ,           T_REG_5__SCAN_IN);
  not   g26( wr_120  ,           X_REG_4__SCAN_IN);
  not   g27( wr_130  ,           CONT_REG_4__SCAN_IN);
  not   g28( wr_101  ,           X_REG_5__SCAN_IN);
  not   g29( wr_113  ,           CONT_REG_5__SCAN_IN);
  not   g30( wr_73   ,           MAR_REG_1__SCAN_IN);
  not   g31( wr_74   ,           MAR_REG_0__SCAN_IN);
  not   g32( wr_217  ,           Y_REG_6__SCAN_IN);
  not   g33( wr_219  ,           T_REG_6__SCAN_IN);
  nor   g34( wr_239  , X_REG_4__SCAN_IN, X_REG_5__SCAN_IN);
  not   g35( wr_72   ,           MAR_REG_2__SCAN_IN);
  not   g36( wr_89   ,           X_REG_6__SCAN_IN);
  not   g37( wr_96   ,           CONT_REG_6__SCAN_IN);
  nor   g38( wr_245  , X_REG_0__SCAN_IN, X_REG_3__SCAN_IN);
  nor   g39( wr_83   , STATO_REG_2__SCAN_IN, STATO_REG_1__SCAN_IN);
  nor   g40( wr_443  , MAR_REG_2__SCAN_IN, MAR_REG_3__SCAN_IN);
  not   g41( wr_230  ,           CONT_REG_7__SCAN_IN);
  nor   g42( wr_431  , STATO_REG_2__SCAN_IN, STATO_REG_0__SCAN_IN);
  nor   g43( wr_500  , MAR_REG_1__SCAN_IN, MAR_REG_3__SCAN_IN);
  not   g44( wr_362  ,           PUNTI_RETTA_REG_0__SCAN_IN);
  not   g45( wr_453  ,           X_REG_7__SCAN_IN);
  not   g46( wr_58   ,           PUNTI_RETTA_REG_7__SCAN_IN);
  not   g47( wr_262  ,           PUNTI_RETTA_REG_6__SCAN_IN);
  not   g48( wr_278  ,           PUNTI_RETTA_REG_5__SCAN_IN);
  not   g49( wr_294  ,           PUNTI_RETTA_REG_4__SCAN_IN);
  not   g50( wr_310  ,           PUNTI_RETTA_REG_3__SCAN_IN);
  not   g51( wr_326  ,           PUNTI_RETTA_REG_2__SCAN_IN);
  not   g52( wr_342  ,           PUNTI_RETTA_REG_1__SCAN_IN);
  not   g53( wr_398  ,           MAR_REG_7__SCAN_IN);
  not   g54( wr_402  ,           MAR_REG_6__SCAN_IN);
  not   g55( wr_403  ,           MAR_REG_5__SCAN_IN);
  not   g56( wr_404  ,           MAR_REG_4__SCAN_IN);
  not   g57( PUNTI_RETTA_7_,           PUNTI_RETTA_REG_7__SCAN_IN);
  not   g58( PUNTI_RETTA_6_,           PUNTI_RETTA_REG_6__SCAN_IN);
  not   g59( PUNTI_RETTA_5_,           PUNTI_RETTA_REG_5__SCAN_IN);
  not   g60( PUNTI_RETTA_4_,           PUNTI_RETTA_REG_4__SCAN_IN);
  not   g61( PUNTI_RETTA_3_,           PUNTI_RETTA_REG_3__SCAN_IN);
  not   g62( PUNTI_RETTA_2_,           PUNTI_RETTA_REG_2__SCAN_IN);
  not   g63( PUNTI_RETTA_1_,           PUNTI_RETTA_REG_1__SCAN_IN);
  not   g64( PUNTI_RETTA_0_,           PUNTI_RETTA_REG_0__SCAN_IN);
  nor   g65( wr_61   , wr_60   , wr_59   );
  nor   g66( wr_90   , wr_60   , wr_82   );
  nor   g67( wr_92   , wr_91   , wr_60   );
  nor   g68( wr_97   , wr_60   , wr_59   );
  not   g69( wr_107  ,           wr_91   );
  nor   g70( wr_155  , STATO_REG_2__SCAN_IN, wr_154  );
  nor   g71( wr_172  , STATO_REG_2__SCAN_IN, wr_171  );
  nor   g72( wr_188  , STATO_REG_2__SCAN_IN, wr_187  );
  nor   g73( wr_138  , STATO_REG_2__SCAN_IN, wr_137  );
  nor   g74( wr_64   , wr_63   , MAR_REG_4__SCAN_IN);
  nor   g75( wr_121  , STATO_REG_2__SCAN_IN, wr_120  );
  nor   g76( wr_102  , STATO_REG_2__SCAN_IN, wr_101  );
  nor   g77( wr_75   , wr_74   , wr_73   );
  not   g78( wr_240  ,           wr_239  );
  nor   g79( wr_216  , STATO_REG_2__SCAN_IN, wr_89   );
  not   g80( wr_246  ,           wr_245  );
  nor   g81( wr_438  , MAR_REG_2__SCAN_IN, wr_63   );
  not   g82( wr_84   ,           wr_83   );
  not   g83( wr_444  ,           wr_443  );
  not   g84( wr_432  ,           wr_431  );
  nor   g85( wr_399  , wr_59   , wr_82   );
  nor   g86( wr_434  , wr_60   , STATO_REG_1__SCAN_IN);
  not   g87( wr_501  ,           wr_500  );
  nor   g88( wr_424  , wr_83   , MAR_REG_0__SCAN_IN);
  nor   g89( wr_488  , wr_74   , MAR_REG_1__SCAN_IN);
  not   g90( wr_93   ,           wr_92   );
  not   g91( wr_98   ,           wr_97   );
  not   g92( wr_104  ,           wr_90   );
  nor   g93( wr_142  , wr_107  , wr_141  );
  nor   g94( wr_159  , wr_107  , wr_158  );
  nor   g95( wr_176  , wr_107  , wr_175  );
  nor   g96( wr_190  , wr_107  , wr_189  );
  nor   g97( wr_125  , wr_107  , wr_124  );
  nor   g98( wr_108  , wr_107  , wr_106  );
  not   g99( wr_65   ,           wr_64   );
  not  g100( wr_76   ,           wr_75   );
  nor  g101( wr_220  , wr_107  , wr_219  );
  nor  g102( wr_241  , wr_240  , X_REG_7__SCAN_IN);
  nor  g103( wr_247  , wr_246  , X_REG_2__SCAN_IN);
  not  g104( wr_62   ,           wr_61   );
  not  g105( wr_439  ,           wr_438  );
  nor  g106( wr_85   , wr_84   , wr_82   );
  nor  g107( wr_445  , wr_444  , MAR_REG_1__SCAN_IN);
  nor  g108( wr_433  , wr_432  , wr_59   );
  nor  g109( wr_417  , wr_83   , wr_75   );
  nor  g110( wr_502  , wr_501  , MAR_REG_2__SCAN_IN);
  nor  g111( wr_510  , wr_107  , wr_60   );
  not  g112( wr_520  ,           wr_399  );
  nor  g113( wr_522  , wr_399  , wr_141  );
  nor  g114( wr_525  , wr_399  , wr_106  );
  nor  g115( wr_528  , wr_399  , wr_175  );
  nor  g116( wr_531  , wr_399  , wr_189  );
  nor  g117( wr_534  , wr_399  , wr_124  );
  nor  g118( wr_537  , wr_399  , wr_219  );
  nor  g119( wr_540  , wr_399  , wr_158  );
  nor  g120( wr_552  , wr_434  , wr_399  );
  nor  g121( wr_94   , wr_93   , wr_90   );
  nor  g122( wr_140  , wr_104  , wr_139  );
  nor  g123( wr_157  , wr_104  , wr_156  );
  nor  g124( wr_165  , wr_98   , wr_164  );
  nor  g125( wr_174  , wr_104  , wr_173  );
  nor  g126( wr_182  , wr_98   , wr_181  );
  nor  g127( wr_186  , wr_104  , wr_185  );
  nor  g128( wr_191  , wr_190  , wr_188  );
  nor  g129( wr_198  , wr_98   , wr_197  );
  nor  g130( wr_123  , wr_104  , wr_122  );
  nor  g131( wr_148  , wr_98   , wr_147  );
  nor  g132( wr_105  , wr_104  , wr_103  );
  nor  g133( wr_131  , wr_98   , wr_130  );
  nor  g134( wr_66   , wr_65   , MAR_REG_5__SCAN_IN);
  nor  g135( wr_114  , wr_98   , wr_113  );
  nor  g136( wr_218  , wr_104  , wr_217  );
  nor  g137( wr_77   , wr_76   , wr_72   );
  nor  g138( wr_99   , wr_98   , wr_96   );
  not  g139( wr_242  ,           wr_241  );
  not  g140( wr_248  ,           wr_247  );
  nor  g141( wr_440  , wr_439  , wr_73   );
  nor  g142( wr_231  , wr_98   , wr_230  );
  not  g143( wr_446  ,           wr_445  );
  nor  g144( wr_435  , wr_434  , wr_433  );
  nor  g145( wr_480  , wr_439  , wr_76   );
  not  g146( wr_511  ,           wr_510  );
  nor  g147( wr_513  , wr_510  , wr_139  );
  nor  g148( wr_515  , wr_510  , wr_173  );
  nor  g149( wr_518  , wr_510  , wr_103  );
  nor  g150( wr_542  , wr_510  , wr_122  );
  nor  g151( wr_544  , wr_510  , wr_185  );
  nor  g152( wr_547  , wr_510  , wr_156  );
  nor  g153( wr_550  , wr_510  , wr_217  );
  not  g154( STATO_REG_2__SCAN_OUT,           wr_552  );
  nor  g155( wr_143  , wr_142  , wr_140  );
  nor  g156( wr_160  , wr_159  , wr_157  );
  nor  g157( wr_163  , wr_94   , wr_154  );
  nor  g158( wr_177  , wr_176  , wr_174  );
  nor  g159( wr_180  , wr_94   , wr_171  );
  not  g160( wr_192  ,           wr_191  );
  nor  g161( wr_196  , wr_94   , wr_187  );
  nor  g162( wr_146  , wr_94   , wr_137  );
  nor  g163( wr_126  , wr_125  , wr_123  );
  nor  g164( wr_129  , wr_94   , wr_120  );
  nor  g165( wr_109  , wr_108  , wr_105  );
  nor  g166( wr_112  , wr_94   , wr_101  );
  not  g167( wr_67   ,           wr_66   );
  nor  g168( wr_95   , wr_94   , wr_89   );
  nor  g169( wr_221  , wr_220  , wr_218  );
  not  g170( wr_78   ,           wr_77   );
  nor  g171( wr_243  , wr_242  , X_REG_6__SCAN_IN);
  not  g172( wr_441  ,           wr_440  );
  not  g173( wr_233  ,           wr_231  );
  nor  g174( wr_447  , wr_446  , wr_74   );
  nor  g175( wr_450  , wr_435  , wr_431  );
  not  g176( wr_454  ,           wr_435  );
  nor  g177( wr_410  , wr_83   , wr_77   );
  nor  g178( wr_436  , wr_435  , STATO_REG_2__SCAN_IN);
  not  g179( wr_161  ,           wr_160  );
  nor  g180( wr_166  , wr_165  , wr_163  );
  not  g181( wr_178  ,           wr_177  );
  nor  g182( wr_183  , wr_182  , wr_180  );
  nor  g183( wr_193  , wr_192  , wr_186  );
  nor  g184( wr_199  , wr_198  , wr_196  );
  not  g185( wr_144  ,           wr_143  );
  nor  g186( wr_149  , wr_148  , wr_146  );
  not  g187( wr_127  ,           wr_126  );
  nor  g188( wr_132  , wr_131  , wr_129  );
  not  g189( wr_110  ,           wr_109  );
  nor  g190( wr_115  , wr_114  , wr_112  );
  nor  g191( wr_68   , wr_67   , MAR_REG_6__SCAN_IN);
  nor  g192( wr_100  , wr_99   , wr_95   );
  not  g193( wr_222  ,           wr_221  );
  not  g194( wr_244  ,           wr_243  );
  nor  g195( wr_442  , wr_441  , MAR_REG_0__SCAN_IN);
  nor  g196( wr_489  , wr_78   , wr_63   );
  not  g197( wr_451  ,           wr_450  );
  nor  g198( wr_455  , wr_454  , wr_453  );
  nor  g199( wr_460  , wr_454  , wr_89   );
  nor  g200( wr_465  , wr_454  , wr_101  );
  nor  g201( wr_470  , wr_454  , wr_120  );
  nor  g202( wr_475  , wr_454  , wr_137  );
  nor  g203( wr_484  , wr_454  , wr_154  );
  nor  g204( wr_495  , wr_454  , wr_171  );
  nor  g205( wr_506  , wr_454  , wr_187  );
  not  g206( wr_437  ,           wr_436  );
  nor  g207( wr_162  , wr_161  , wr_155  );
  nor  g208( wr_179  , wr_178  , wr_172  );
  not  g209( wr_194  ,           wr_193  );
  not  g210( wr_203  ,           wr_183  );
  not  g211( wr_169  ,           wr_166  );
  nor  g212( wr_145  , wr_144  , wr_138  );
  not  g213( wr_152  ,           wr_149  );
  nor  g214( wr_128  , wr_127  , wr_121  );
  not  g215( wr_135  ,           wr_132  );
  nor  g216( wr_111  , wr_110  , wr_102  );
  not  g217( wr_118  ,           wr_115  );
  not  g218( wr_69   ,           wr_68   );
  nor  g219( wr_223  , wr_222  , wr_216  );
  not  g220( wr_224  ,           wr_100  );
  nor  g221( wr_249  , wr_248  , wr_244  );
  not  g222( wr_358  ,           wr_199  );
  nor  g223( wr_448  , wr_447  , wr_442  );
  nor  g224( wr_195  , wr_194  , wr_61   );
  not  g225( wr_202  ,           wr_179  );
  not  g226( wr_168  ,           wr_162  );
  nor  g227( wr_184  , wr_183  , wr_179  );
  not  g228( wr_151  ,           wr_145  );
  nor  g229( wr_167  , wr_166  , wr_162  );
  not  g230( wr_134  ,           wr_128  );
  nor  g231( wr_150  , wr_149  , wr_145  );
  not  g232( wr_117  ,           wr_111  );
  nor  g233( wr_133  , wr_132  , wr_128  );
  nor  g234( wr_70   , wr_69   , MAR_REG_7__SCAN_IN);
  nor  g235( wr_116  , wr_115  , wr_111  );
  not  g236( wr_264  ,           wr_223  );
  nor  g237( wr_266  , wr_223  , wr_224  );
  nor  g238( wr_281  , wr_118  , wr_111  );
  nor  g239( wr_297  , wr_135  , wr_128  );
  nor  g240( wr_313  , wr_152  , wr_145  );
  nor  g241( wr_329  , wr_169  , wr_162  );
  not  g242( wr_250  ,           wr_249  );
  nor  g243( wr_344  , wr_203  , wr_179  );
  not  g244( wr_479  ,           wr_448  );
  nor  g245( wr_449  , wr_448  , wr_437  );
  nor  g246( wr_512  , wr_511  , wr_448  );
  nor  g247( wr_200  , wr_199  , wr_195  );
  nor  g248( wr_204  , wr_203  , wr_202  );
  nor  g249( wr_170  , wr_169  , wr_168  );
  nor  g250( wr_153  , wr_152  , wr_151  );
  nor  g251( wr_136  , wr_135  , wr_134  );
  nor  g252( wr_119  , wr_118  , wr_117  );
  not  g253( wr_71   ,           wr_70   );
  nor  g254( wr_265  , wr_264  , wr_100  );
  nor  g255( wr_280  , wr_115  , wr_117  );
  nor  g256( wr_296  , wr_132  , wr_134  );
  nor  g257( wr_312  , wr_149  , wr_151  );
  nor  g258( wr_328  , wr_166  , wr_168  );
  nor  g259( wr_345  , wr_183  , wr_202  );
  nor  g260( wr_251  , wr_250  , wr_171  );
  not  g261( wr_356  ,           wr_195  );
  nor  g262( wr_359  , wr_358  , wr_195  );
  nor  g263( wr_481  , wr_480  , wr_479  );
  nor  g264( wr_490  , wr_489  , wr_479  );
  nor  g265( wr_514  , wr_513  , wr_512  );
  nor  g266( wr_519  , wr_518  , wr_512  );
  nor  g267( wr_543  , wr_542  , wr_512  );
  nor  g268( wr_551  , wr_550  , wr_512  );
  not  g269( wr_201  ,           wr_200  );
  nor  g270( wr_79   , wr_78   , wr_71   );
  nor  g271( wr_267  , wr_266  , wr_265  );
  nor  g272( wr_282  , wr_281  , wr_280  );
  nor  g273( wr_298  , wr_297  , wr_296  );
  nor  g274( wr_314  , wr_313  , wr_312  );
  nor  g275( wr_330  , wr_329  , wr_328  );
  nor  g276( wr_346  , wr_345  , wr_344  );
  not  g277( wr_252  ,           wr_251  );
  nor  g278( wr_357  , wr_199  , wr_356  );
  not  g279( wr_491  ,           wr_490  );
  not  g280( wr_499  ,           wr_481  );
  nor  g281( wr_482  , wr_481  , wr_437  );
  nor  g282( wr_548  , wr_511  , wr_481  );
  not  g283( Y_REG_3__SCAN_OUT,           wr_514  );
  not  g284( Y_REG_5__SCAN_OUT,           wr_519  );
  not  g285( Y_REG_4__SCAN_OUT,           wr_543  );
  not  g286( Y_REG_6__SCAN_OUT,           wr_551  );
  nor  g287( wr_205  , wr_204  , wr_201  );
  not  g288( wr_80   ,           wr_79   );
  not  g289( wr_269  ,           wr_267  );
  not  g290( wr_285  ,           wr_282  );
  not  g291( wr_301  ,           wr_298  );
  not  g292( wr_317  ,           wr_314  );
  not  g293( wr_333  ,           wr_330  );
  nor  g294( wr_368  , wr_79   , wr_62   );
  not  g295( wr_348  ,           wr_346  );
  nor  g296( wr_347  , wr_346  , wr_200  );
  nor  g297( wr_360  , wr_359  , wr_357  );
  nor  g298( wr_553  , wr_79   , STATO_REG_0__SCAN_IN);
  nor  g299( wr_492  , wr_491  , wr_488  );
  nor  g300( wr_503  , wr_502  , wr_499  );
  nor  g301( wr_549  , wr_548  , wr_547  );
  nor  g302( wr_206  , wr_205  , wr_184  );
  nor  g303( wr_81   , wr_80   , wr_62   );
  not  g304( wr_369  ,           wr_368  );
  nor  g305( wr_400  , wr_399  , wr_368  );
  nor  g306( wr_349  , wr_348  , wr_201  );
  nor  g307( wr_505  , wr_451  , wr_360  );
  nor  g308( wr_554  , wr_553  , wr_431  );
  nor  g309( wr_493  , wr_492  , wr_437  );
  nor  g310( wr_504  , wr_503  , wr_437  );
  nor  g311( wr_516  , wr_511  , wr_492  );
  nor  g312( wr_530  , wr_520  , wr_360  );
  nor  g313( wr_545  , wr_511  , wr_503  );
  not  g314( Y_REG_2__SCAN_OUT,           wr_549  );
  nor  g315( wr_207  , wr_206  , wr_170  );
  nor  g316( wr_86   , wr_85   , wr_81   );
  not  g317( wr_332  ,           wr_206  );
  nor  g318( wr_331  , wr_330  , wr_206  );
  nor  g319( wr_370  , wr_252  , wr_369  );
  nor  g320( wr_405  , wr_400  , wr_83   );
  nor  g321( wr_350  , wr_349  , wr_347  );
  nor  g322( wr_557  , wr_83   , wr_81   );
  not  g323( wr_401  ,           wr_400  );
  nor  g324( wr_411  , wr_410  , wr_400  );
  nor  g325( wr_418  , wr_417  , wr_400  );
  nor  g326( wr_425  , wr_424  , wr_400  );
  nor  g327( wr_507  , wr_506  , wr_505  );
  nor  g328( wr_555  , wr_554  , wr_59   );
  nor  g329( wr_517  , wr_516  , wr_515  );
  nor  g330( wr_532  , wr_531  , wr_530  );
  nor  g331( wr_546  , wr_545  , wr_544  );
  nor  g332( wr_208  , wr_207  , wr_167  );
  nor  g333( wr_237  , wr_86   , wr_60   );
  nor  g334( wr_334  , wr_333  , wr_332  );
  not  g335( wr_87   ,           wr_86   );
  not  g336( wr_372  ,           wr_370  );
  not  g337( wr_406  ,           wr_405  );
  nor  g338( wr_494  , wr_451  , wr_350  );
  not  g339( wr_558  ,           wr_557  );
  nor  g340( wr_371  , wr_370  , wr_230  );
  nor  g341( wr_377  , wr_370  , wr_96   );
  nor  g342( wr_380  , wr_370  , wr_113  );
  nor  g343( wr_383  , wr_370  , wr_130  );
  nor  g344( wr_386  , wr_370  , wr_147  );
  nor  g345( wr_389  , wr_370  , wr_164  );
  nor  g346( wr_392  , wr_370  , wr_181  );
  nor  g347( wr_395  , wr_370  , wr_197  );
  nor  g348( wr_412  , wr_411  , wr_63   );
  nor  g349( wr_419  , wr_418  , wr_72   );
  nor  g350( wr_426  , wr_425  , wr_73   );
  nor  g351( wr_428  , wr_401  , wr_74   );
  not  g352( wr_508  ,           wr_507  );
  nor  g353( wr_527  , wr_520  , wr_350  );
  nor  g354( wr_556  , wr_555  , wr_90   );
  nor  g355( MAR_REG_7__SCAN_OUT, wr_401  , wr_398  );
  nor  g356( MAR_REG_6__SCAN_OUT, wr_401  , wr_402  );
  nor  g357( MAR_REG_5__SCAN_OUT, wr_401  , wr_403  );
  nor  g358( MAR_REG_4__SCAN_OUT, wr_401  , wr_404  );
  not  g359( Y_REG_1__SCAN_OUT,           wr_517  );
  not  g360( T_REG_0__SCAN_OUT,           wr_532  );
  not  g361( Y_REG_0__SCAN_OUT,           wr_546  );
  nor  g362( wr_209  , wr_208  , wr_153  );
  not  g363( wr_316  ,           wr_208  );
  not  g364( wr_238  ,           wr_237  );
  nor  g365( wr_315  , wr_314  , wr_208  );
  nor  g366( wr_335  , wr_334  , wr_331  );
  nor  g367( wr_363  , wr_87   , wr_362  );
  nor  g368( wr_373  , wr_372  , wr_60   );
  nor  g369( wr_407  , wr_406  , MAR_REG_3__SCAN_IN);
  nor  g370( wr_414  , wr_406  , MAR_REG_2__SCAN_IN);
  nor  g371( wr_421  , wr_406  , wr_74   );
  nor  g372( wr_496  , wr_495  , wr_494  );
  nor  g373( wr_559  , wr_558  , wr_431  );
  nor  g374( wr_88   , wr_87   , wr_58   );
  nor  g375( wr_263  , wr_87   , wr_262  );
  nor  g376( wr_279  , wr_87   , wr_278  );
  nor  g377( wr_295  , wr_87   , wr_294  );
  nor  g378( wr_311  , wr_87   , wr_310  );
  nor  g379( wr_327  , wr_87   , wr_326  );
  nor  g380( wr_343  , wr_87   , wr_342  );
  nor  g381( wr_429  , wr_406  , MAR_REG_0__SCAN_IN);
  nor  g382( wr_509  , wr_508  , wr_504  );
  nor  g383( wr_529  , wr_528  , wr_527  );
  not  g384( STATO_REG_1__SCAN_OUT,           wr_556  );
  nor  g385( wr_210  , wr_209  , wr_150  );
  nor  g386( wr_318  , wr_317  , wr_316  );
  nor  g387( wr_253  , wr_252  , wr_238  );
  nor  g388( wr_256  , wr_251  , wr_238  );
  not  g389( wr_336  ,           wr_335  );
  not  g390( wr_374  ,           wr_373  );
  not  g391( wr_408  ,           wr_407  );
  not  g392( wr_415  ,           wr_414  );
  not  g393( wr_422  ,           wr_421  );
  not  g394( wr_497  ,           wr_496  );
  not  g395( wr_560  ,           wr_559  );
  nor  g396( wr_430  , wr_429  , wr_428  );
  not  g397( X_REG_0__SCAN_OUT,           wr_509  );
  not  g398( T_REG_1__SCAN_OUT,           wr_529  );
  nor  g399( wr_211  , wr_210  , wr_136  );
  not  g400( wr_300  ,           wr_210  );
  nor  g401( wr_299  , wr_298  , wr_210  );
  nor  g402( wr_319  , wr_318  , wr_315  );
  not  g403( wr_254  ,           wr_253  );
  not  g404( wr_257  ,           wr_256  );
  nor  g405( wr_483  , wr_451  , wr_336  );
  nor  g406( wr_390  , wr_374  , wr_336  );
  nor  g407( wr_393  , wr_374  , wr_350  );
  nor  g408( wr_396  , wr_374  , wr_360  );
  nor  g409( wr_409  , wr_408  , wr_78   );
  nor  g410( wr_416  , wr_415  , wr_76   );
  nor  g411( wr_423  , wr_422  , MAR_REG_1__SCAN_IN);
  nor  g412( wr_539  , wr_520  , wr_336  );
  nor  g413( wr_498  , wr_497  , wr_493  );
  nor  g414( wr_561  , wr_560  , wr_91   );
  not  g415( MAR_REG_0__SCAN_OUT,           wr_430  );
  nor  g416( wr_212  , wr_211  , wr_133  );
  nor  g417( wr_302  , wr_301  , wr_300  );
  not  g418( wr_320  ,           wr_319  );
  nor  g419( wr_258  , wr_257  , wr_230  );
  nor  g420( wr_274  , wr_257  , wr_96   );
  nor  g421( wr_290  , wr_257  , wr_113  );
  nor  g422( wr_306  , wr_257  , wr_130  );
  nor  g423( wr_322  , wr_257  , wr_147  );
  nor  g424( wr_337  , wr_336  , wr_254  );
  nor  g425( wr_338  , wr_257  , wr_164  );
  nor  g426( wr_351  , wr_350  , wr_254  );
  nor  g427( wr_352  , wr_257  , wr_181  );
  nor  g428( wr_364  , wr_257  , wr_197  );
  nor  g429( wr_485  , wr_484  , wr_483  );
  nor  g430( wr_361  , wr_360  , wr_254  );
  nor  g431( wr_391  , wr_390  , wr_389  );
  nor  g432( wr_394  , wr_393  , wr_392  );
  nor  g433( wr_397  , wr_396  , wr_395  );
  nor  g434( wr_413  , wr_412  , wr_409  );
  nor  g435( wr_420  , wr_419  , wr_416  );
  nor  g436( wr_427  , wr_426  , wr_423  );
  nor  g437( wr_541  , wr_540  , wr_539  );
  not  g438( X_REG_1__SCAN_OUT,           wr_498  );
  not  g439( STATO_REG_0__SCAN_OUT,           wr_561  );
  nor  g440( wr_213  , wr_212  , wr_119  );
  not  g441( wr_284  ,           wr_212  );
  nor  g442( wr_283  , wr_282  , wr_212  );
  nor  g443( wr_303  , wr_302  , wr_299  );
  nor  g444( wr_321  , wr_320  , wr_254  );
  nor  g445( wr_474  , wr_451  , wr_320  );
  nor  g446( wr_339  , wr_338  , wr_337  );
  nor  g447( wr_353  , wr_352  , wr_351  );
  nor  g448( wr_365  , wr_364  , wr_363  );
  nor  g449( wr_387  , wr_374  , wr_320  );
  not  g450( wr_486  ,           wr_485  );
  nor  g451( wr_521  , wr_520  , wr_320  );
  not  g452( CONT_REG_2__SCAN_OUT,           wr_391  );
  not  g453( CONT_REG_1__SCAN_OUT,           wr_394  );
  not  g454( CONT_REG_0__SCAN_OUT,           wr_397  );
  not  g455( MAR_REG_3__SCAN_OUT,           wr_413  );
  not  g456( MAR_REG_2__SCAN_OUT,           wr_420  );
  not  g457( MAR_REG_1__SCAN_OUT,           wr_427  );
  not  g458( T_REG_2__SCAN_OUT,           wr_541  );
  nor  g459( wr_214  , wr_213  , wr_116  );
  nor  g460( wr_286  , wr_285  , wr_284  );
  not  g461( wr_304  ,           wr_303  );
  nor  g462( wr_323  , wr_322  , wr_321  );
  nor  g463( wr_476  , wr_475  , wr_474  );
  not  g464( wr_340  ,           wr_339  );
  not  g465( wr_354  ,           wr_353  );
  not  g466( wr_366  ,           wr_365  );
  nor  g467( wr_388  , wr_387  , wr_386  );
  nor  g468( wr_487  , wr_486  , wr_482  );
  nor  g469( wr_523  , wr_522  , wr_521  );
  not  g470( wr_225  ,           wr_214  );
  nor  g471( wr_215  , wr_214  , wr_100  );
  nor  g472( wr_268  , wr_267  , wr_214  );
  nor  g473( wr_287  , wr_286  , wr_283  );
  nor  g474( wr_305  , wr_304  , wr_254  );
  nor  g475( wr_469  , wr_451  , wr_304  );
  not  g476( wr_324  ,           wr_323  );
  nor  g477( wr_384  , wr_374  , wr_304  );
  not  g478( wr_477  ,           wr_476  );
  nor  g479( wr_533  , wr_520  , wr_304  );
  nor  g480( wr_341  , wr_340  , wr_327  );
  nor  g481( wr_355  , wr_354  , wr_343  );
  nor  g482( wr_367  , wr_366  , wr_361  );
  not  g483( CONT_REG_3__SCAN_OUT,           wr_388  );
  not  g484( X_REG_2__SCAN_OUT,           wr_487  );
  not  g485( T_REG_3__SCAN_OUT,           wr_523  );
  nor  g486( wr_226  , wr_225  , wr_224  );
  nor  g487( wr_270  , wr_269  , wr_225  );
  not  g488( wr_288  ,           wr_287  );
  nor  g489( wr_307  , wr_306  , wr_305  );
  nor  g490( wr_471  , wr_470  , wr_469  );
  nor  g491( wr_325  , wr_324  , wr_311  );
  nor  g492( wr_385  , wr_384  , wr_383  );
  nor  g493( wr_478  , wr_477  , wr_449  );
  nor  g494( wr_535  , wr_534  , wr_533  );
  not  g495( PUNTI_RETTA_REG_2__SCAN_OUT,           wr_341  );
  not  g496( PUNTI_RETTA_REG_1__SCAN_OUT,           wr_355  );
  not  g497( PUNTI_RETTA_REG_0__SCAN_OUT,           wr_367  );
  nor  g498( wr_227  , wr_226  , wr_223  );
  nor  g499( wr_271  , wr_270  , wr_268  );
  nor  g500( wr_289  , wr_288  , wr_254  );
  nor  g501( wr_464  , wr_451  , wr_288  );
  not  g502( wr_308  ,           wr_307  );
  nor  g503( wr_381  , wr_374  , wr_288  );
  not  g504( wr_472  ,           wr_471  );
  nor  g505( wr_524  , wr_520  , wr_288  );
  not  g506( PUNTI_RETTA_REG_3__SCAN_OUT,           wr_325  );
  not  g507( CONT_REG_4__SCAN_OUT,           wr_385  );
  not  g508( X_REG_3__SCAN_OUT,           wr_478  );
  not  g509( T_REG_4__SCAN_OUT,           wr_535  );
  nor  g510( wr_228  , wr_227  , wr_215  );
  not  g511( wr_272  ,           wr_271  );
  nor  g512( wr_291  , wr_290  , wr_289  );
  nor  g513( wr_466  , wr_465  , wr_464  );
  nor  g514( wr_309  , wr_308  , wr_295  );
  nor  g515( wr_382  , wr_381  , wr_380  );
  nor  g516( wr_473  , wr_472  , wr_449  );
  nor  g517( wr_526  , wr_525  , wr_524  );
  not  g518( wr_229  ,           wr_228  );
  nor  g519( wr_234  , wr_233  , wr_228  );
  nor  g520( wr_273  , wr_272  , wr_254  );
  nor  g521( wr_459  , wr_451  , wr_272  );
  not  g522( wr_292  ,           wr_291  );
  nor  g523( wr_378  , wr_374  , wr_272  );
  not  g524( wr_467  ,           wr_466  );
  nor  g525( wr_536  , wr_520  , wr_272  );
  not  g526( PUNTI_RETTA_REG_4__SCAN_OUT,           wr_309  );
  not  g527( CONT_REG_5__SCAN_OUT,           wr_382  );
  not  g528( X_REG_4__SCAN_OUT,           wr_473  );
  not  g529( T_REG_5__SCAN_OUT,           wr_526  );
  nor  g530( wr_232  , wr_231  , wr_229  );
  nor  g531( wr_275  , wr_274  , wr_273  );
  nor  g532( wr_461  , wr_460  , wr_459  );
  nor  g533( wr_293  , wr_292  , wr_279  );
  nor  g534( wr_379  , wr_378  , wr_377  );
  nor  g535( wr_468  , wr_467  , wr_449  );
  nor  g536( wr_538  , wr_537  , wr_536  );
  nor  g537( wr_235  , wr_234  , wr_232  );
  not  g538( wr_276  ,           wr_275  );
  not  g539( wr_462  ,           wr_461  );
  not  g540( PUNTI_RETTA_REG_5__SCAN_OUT,           wr_293  );
  not  g541( CONT_REG_6__SCAN_OUT,           wr_379  );
  not  g542( X_REG_5__SCAN_OUT,           wr_468  );
  not  g543( T_REG_6__SCAN_OUT,           wr_538  );
  not  g544( wr_236  ,           wr_235  );
  nor  g545( wr_277  , wr_276  , wr_263  );
  nor  g546( wr_463  , wr_462  , wr_449  );
  nor  g547( wr_255  , wr_254  , wr_236  );
  nor  g548( wr_452  , wr_451  , wr_236  );
  nor  g549( wr_375  , wr_374  , wr_236  );
  not  g550( PUNTI_RETTA_REG_6__SCAN_OUT,           wr_277  );
  not  g551( X_REG_6__SCAN_OUT,           wr_463  );
  nor  g552( wr_259  , wr_258  , wr_255  );
  nor  g553( wr_456  , wr_455  , wr_452  );
  nor  g554( wr_376  , wr_375  , wr_371  );
  not  g555( wr_260  ,           wr_259  );
  not  g556( wr_457  ,           wr_456  );
  not  g557( CONT_REG_7__SCAN_OUT,           wr_376  );
  nor  g558( wr_261  , wr_260  , wr_88   );
  nor  g559( wr_458  , wr_457  , wr_449  );
  not  g560( PUNTI_RETTA_REG_7__SCAN_OUT,           wr_261  );
  not  g561( X_REG_7__SCAN_OUT,           wr_458  );

endmodule
