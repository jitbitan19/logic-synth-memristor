// NOR_NOT mapped module c5315

module c5315 (
  input  G1      ,
  input  G4      ,
  input  G11     ,
  input  G14     ,
  input  G17     ,
  input  G20     ,
  input  G23     ,
  input  G24     ,
  input  G25     ,
  input  G26     ,
  input  G27     ,
  input  G31     ,
  input  G34     ,
  input  G37     ,
  input  G40     ,
  input  G43     ,
  input  G46     ,
  input  G49     ,
  input  G52     ,
  input  G53     ,
  input  G54     ,
  input  G61     ,
  input  G64     ,
  input  G67     ,
  input  G70     ,
  input  G73     ,
  input  G76     ,
  input  G79     ,
  input  G80     ,
  input  G81     ,
  input  G82     ,
  input  G83     ,
  input  G86     ,
  input  G87     ,
  input  G88     ,
  input  G91     ,
  input  G94     ,
  input  G97     ,
  input  G100    ,
  input  G103    ,
  input  G106    ,
  input  G109    ,
  input  G112    ,
  input  G113    ,
  input  G114    ,
  input  G115    ,
  input  G116    ,
  input  G117    ,
  input  G118    ,
  input  G119    ,
  input  G120    ,
  input  G121    ,
  input  G122    ,
  input  G123    ,
  input  G126    ,
  input  G127    ,
  input  G128    ,
  input  G129    ,
  input  G130    ,
  input  G131    ,
  input  G132    ,
  input  G135    ,
  input  G136    ,
  input  G137    ,
  input  G140    ,
  input  G141    ,
  input  G145    ,
  input  G146    ,
  input  G149    ,
  input  G152    ,
  input  G155    ,
  input  G158    ,
  input  G161    ,
  input  G164    ,
  input  G167    ,
  input  G170    ,
  input  G173    ,
  input  G176    ,
  input  G179    ,
  input  G182    ,
  input  G185    ,
  input  G188    ,
  input  G191    ,
  input  G194    ,
  input  G197    ,
  input  G200    ,
  input  G203    ,
  input  G206    ,
  input  G209    ,
  input  G210    ,
  input  G217    ,
  input  G218    ,
  input  G225    ,
  input  G226    ,
  input  G233    ,
  input  G234    ,
  input  G241    ,
  input  G242    ,
  input  G245    ,
  input  G248    ,
  input  G251    ,
  input  G254    ,
  input  G257    ,
  input  G264    ,
  input  G265    ,
  input  G272    ,
  input  G273    ,
  input  G280    ,
  input  G281    ,
  input  G288    ,
  input  G289    ,
  input  G292    ,
  input  G293    ,
  input  G299    ,
  input  G302    ,
  input  G307    ,
  input  G308    ,
  input  G315    ,
  input  G316    ,
  input  G323    ,
  input  G324    ,
  input  G331    ,
  input  G332    ,
  input  G335    ,
  input  G338    ,
  input  G341    ,
  input  G348    ,
  input  G351    ,
  input  G358    ,
  input  G361    ,
  input  G366    ,
  input  G369    ,
  input  G372    ,
  input  G373    ,
  input  G374    ,
  input  G386    ,
  input  G389    ,
  input  G400    ,
  input  G411    ,
  input  G422    ,
  input  G435    ,
  input  G446    ,
  input  G457    ,
  input  G468    ,
  input  G479    ,
  input  G490    ,
  input  G503    ,
  input  G514    ,
  input  G523    ,
  input  G534    ,
  input  G545    ,
  input  G549    ,
  input  G552    ,
  input  G556    ,
  input  G559    ,
  input  G562    ,
  input  G1497   ,
  input  G1689   ,
  input  G1690   ,
  input  G1691   ,
  input  G1694   ,
  input  G2174   ,
  input  G2358   ,
  input  G2824   ,
  input  G3173   ,
  input  G3546   ,
  input  G3548   ,
  input  G3550   ,
  input  G3552   ,
  input  G3717   ,
  input  G3724   ,
  input  G4087   ,
  input  G4088   ,
  input  G4089   ,
  input  G4090   ,
  input  G4091   ,
  input  G4092   ,
  input  G4115   ,
  output G144    ,
  output G298    ,
  output G973    ,
  output G594    ,
  output G599    ,
  output G600    ,
  output G601    ,
  output G602    ,
  output G603    ,
  output G604    ,
  output G611    ,
  output G612    ,
  output G810    ,
  output G848    ,
  output G849    ,
  output G850    ,
  output G851    ,
  output G634    ,
  output G815    ,
  output G845    ,
  output G847    ,
  output G926    ,
  output G923    ,
  output G921    ,
  output G892    ,
  output G887    ,
  output G606    ,
  output G656    ,
  output G809    ,
  output G993    ,
  output G978    ,
  output G949    ,
  output G939    ,
  output G889    ,
  output G593    ,
  output G636    ,
  output G704    ,
  output G717    ,
  output G820    ,
  output G639    ,
  output G673    ,
  output G707    ,
  output G715    ,
  output G598    ,
  output G610    ,
  output G588    ,
  output G615    ,
  output G626    ,
  output G632    ,
  output G1002   ,
  output G1004   ,
  output G591    ,
  output G618    ,
  output G621    ,
  output G629    ,
  output G822    ,
  output G838    ,
  output G861    ,
  output G623    ,
  output G722    ,
  output G832    ,
  output G834    ,
  output G836    ,
  output G859    ,
  output G871    ,
  output G873    ,
  output G875    ,
  output G877    ,
  output G998    ,
  output G1000   ,
  output G575    ,
  output G585    ,
  output G661    ,
  output G693    ,
  output G747    ,
  output G752    ,
  output G757    ,
  output G762    ,
  output G787    ,
  output G792    ,
  output G797    ,
  output G802    ,
  output G642    ,
  output G664    ,
  output G667    ,
  output G670    ,
  output G676    ,
  output G696    ,
  output G699    ,
  output G702    ,
  output G818    ,
  output G813    ,
  output G824    ,
  output G826    ,
  output G828    ,
  output G830    ,
  output G854    ,
  output G863    ,
  output G865    ,
  output G867    ,
  output G869    ,
  output G712    ,
  output G727    ,
  output G732    ,
  output G737    ,
  output G742    ,
  output G772    ,
  output G777    ,
  output G782    ,
  output G645    ,
  output G648    ,
  output G651    ,
  output G654    ,
  output G679    ,
  output G682    ,
  output G685    ,
  output G688    ,
  output G843    ,
  output G882    ,
  output G767    ,
  output G807    ,
  output G658    ,
  output G690    );

  wire wr_124;
  wire wr_125;
  wire wr_126;
  wire wr_127;
  wire wr_128;
  wire wr_129;
  wire wr_130;
  wire wr_131;
  wire wr_132;
  wire wr_133;
  wire wr_134;
  wire wr_135;
  wire wr_136;
  wire wr_137;
  wire wr_138;
  wire wr_139;
  wire wr_140;
  wire wr_141;
  wire wr_142;
  wire wr_143;
  wire wr_144;
  wire wr_145;
  wire wr_146;
  wire wr_147;
  wire wr_148;
  wire wr_149;
  wire wr_150;
  wire wr_151;
  wire wr_152;
  wire wr_153;
  wire wr_154;
  wire wr_155;
  wire wr_156;
  wire wr_157;
  wire wr_158;
  wire wr_159;
  wire wr_160;
  wire wr_161;
  wire wr_162;
  wire wr_163;
  wire wr_164;
  wire wr_165;
  wire wr_166;
  wire wr_167;
  wire wr_168;
  wire wr_169;
  wire wr_170;
  wire wr_171;
  wire wr_172;
  wire wr_173;
  wire wr_174;
  wire wr_175;
  wire wr_176;
  wire wr_177;
  wire wr_178;
  wire wr_179;
  wire wr_180;
  wire wr_181;
  wire wr_182;
  wire wr_183;
  wire wr_184;
  wire wr_185;
  wire wr_186;
  wire wr_187;
  wire wr_188;
  wire wr_189;
  wire wr_190;
  wire wr_191;
  wire wr_192;
  wire wr_193;
  wire wr_194;
  wire wr_195;
  wire wr_196;
  wire wr_197;
  wire wr_198;
  wire wr_199;
  wire wr_200;
  wire wr_201;
  wire wr_202;
  wire wr_203;
  wire wr_204;
  wire wr_205;
  wire wr_206;
  wire wr_207;
  wire wr_208;
  wire wr_209;
  wire wr_210;
  wire wr_211;
  wire wr_212;
  wire wr_213;
  wire wr_214;
  wire wr_215;
  wire wr_216;
  wire wr_217;
  wire wr_218;
  wire wr_219;
  wire wr_220;
  wire wr_221;
  wire wr_222;
  wire wr_223;
  wire wr_224;
  wire wr_225;
  wire wr_226;
  wire wr_227;
  wire wr_228;
  wire wr_229;
  wire wr_230;
  wire wr_231;
  wire wr_232;
  wire wr_233;
  wire wr_234;
  wire wr_235;
  wire wr_236;
  wire wr_237;
  wire wr_238;
  wire wr_239;
  wire wr_240;
  wire wr_241;
  wire wr_242;
  wire wr_243;
  wire wr_244;
  wire wr_245;
  wire wr_246;
  wire wr_247;
  wire wr_248;
  wire wr_249;
  wire wr_250;
  wire wr_251;
  wire wr_252;
  wire wr_253;
  wire wr_254;
  wire wr_255;
  wire wr_256;
  wire wr_257;
  wire wr_258;
  wire wr_259;
  wire wr_260;
  wire wr_261;
  wire wr_262;
  wire wr_263;
  wire wr_264;
  wire wr_265;
  wire wr_266;
  wire wr_267;
  wire wr_268;
  wire wr_269;
  wire wr_270;
  wire wr_271;
  wire wr_272;
  wire wr_273;
  wire wr_274;
  wire wr_275;
  wire wr_276;
  wire wr_277;
  wire wr_278;
  wire wr_279;
  wire wr_280;
  wire wr_281;
  wire wr_282;
  wire wr_283;
  wire wr_284;
  wire wr_285;
  wire wr_286;
  wire wr_287;
  wire wr_288;
  wire wr_289;
  wire wr_290;
  wire wr_291;
  wire wr_292;
  wire wr_293;
  wire wr_294;
  wire wr_295;
  wire wr_296;
  wire wr_297;
  wire wr_298;
  wire wr_299;
  wire wr_300;
  wire wr_301;
  wire wr_302;
  wire wr_303;
  wire wr_304;
  wire wr_305;
  wire wr_306;
  wire wr_307;
  wire wr_308;
  wire wr_309;
  wire wr_310;
  wire wr_311;
  wire wr_312;
  wire wr_313;
  wire wr_314;
  wire wr_315;
  wire wr_316;
  wire wr_317;
  wire wr_318;
  wire wr_319;
  wire wr_320;
  wire wr_321;
  wire wr_322;
  wire wr_323;
  wire wr_324;
  wire wr_325;
  wire wr_326;
  wire wr_327;
  wire wr_328;
  wire wr_329;
  wire wr_330;
  wire wr_331;
  wire wr_332;
  wire wr_333;
  wire wr_334;
  wire wr_335;
  wire wr_336;
  wire wr_337;
  wire wr_338;
  wire wr_339;
  wire wr_340;
  wire wr_341;
  wire wr_342;
  wire wr_343;
  wire wr_344;
  wire wr_345;
  wire wr_346;
  wire wr_347;
  wire wr_348;
  wire wr_349;
  wire wr_350;
  wire wr_351;
  wire wr_352;
  wire wr_353;
  wire wr_354;
  wire wr_355;
  wire wr_356;
  wire wr_357;
  wire wr_358;
  wire wr_359;
  wire wr_360;
  wire wr_361;
  wire wr_362;
  wire wr_363;
  wire wr_364;
  wire wr_365;
  wire wr_366;
  wire wr_367;
  wire wr_368;
  wire wr_369;
  wire wr_370;
  wire wr_371;
  wire wr_372;
  wire wr_373;
  wire wr_374;
  wire wr_375;
  wire wr_376;
  wire wr_377;
  wire wr_378;
  wire wr_379;
  wire wr_380;
  wire wr_381;
  wire wr_382;
  wire wr_383;
  wire wr_384;
  wire wr_385;
  wire wr_386;
  wire wr_387;
  wire wr_388;
  wire wr_389;
  wire wr_390;
  wire wr_391;
  wire wr_392;
  wire wr_393;
  wire wr_394;
  wire wr_395;
  wire wr_396;
  wire wr_397;
  wire wr_398;
  wire wr_399;
  wire wr_400;
  wire wr_401;
  wire wr_402;
  wire wr_403;
  wire wr_404;
  wire wr_405;
  wire wr_406;
  wire wr_407;
  wire wr_408;
  wire wr_409;
  wire wr_410;
  wire wr_411;
  wire wr_412;
  wire wr_413;
  wire wr_414;
  wire wr_415;
  wire wr_416;
  wire wr_417;
  wire wr_418;
  wire wr_419;
  wire wr_420;
  wire wr_421;
  wire wr_422;
  wire wr_423;
  wire wr_424;
  wire wr_425;
  wire wr_426;
  wire wr_427;
  wire wr_428;
  wire wr_429;
  wire wr_430;
  wire wr_431;
  wire wr_432;
  wire wr_433;
  wire wr_434;
  wire wr_435;
  wire wr_436;
  wire wr_437;
  wire wr_438;
  wire wr_439;
  wire wr_440;
  wire wr_441;
  wire wr_442;
  wire wr_443;
  wire wr_444;
  wire wr_445;
  wire wr_446;
  wire wr_447;
  wire wr_448;
  wire wr_449;
  wire wr_450;
  wire wr_451;
  wire wr_452;
  wire wr_453;
  wire wr_454;
  wire wr_455;
  wire wr_456;
  wire wr_457;
  wire wr_458;
  wire wr_459;
  wire wr_460;
  wire wr_461;
  wire wr_462;
  wire wr_463;
  wire wr_464;
  wire wr_465;
  wire wr_466;
  wire wr_467;
  wire wr_468;
  wire wr_469;
  wire wr_470;
  wire wr_471;
  wire wr_472;
  wire wr_473;
  wire wr_474;
  wire wr_475;
  wire wr_476;
  wire wr_477;
  wire wr_478;
  wire wr_479;
  wire wr_480;
  wire wr_481;
  wire wr_482;
  wire wr_483;
  wire wr_484;
  wire wr_485;
  wire wr_486;
  wire wr_487;
  wire wr_488;
  wire wr_489;
  wire wr_490;
  wire wr_491;
  wire wr_492;
  wire wr_493;
  wire wr_494;
  wire wr_495;
  wire wr_496;
  wire wr_497;
  wire wr_498;
  wire wr_499;
  wire wr_500;
  wire wr_501;
  wire wr_502;
  wire wr_503;
  wire wr_504;
  wire wr_505;
  wire wr_506;
  wire wr_507;
  wire wr_508;
  wire wr_509;
  wire wr_510;
  wire wr_511;
  wire wr_512;
  wire wr_513;
  wire wr_514;
  wire wr_515;
  wire wr_516;
  wire wr_517;
  wire wr_518;
  wire wr_519;
  wire wr_520;
  wire wr_521;
  wire wr_522;
  wire wr_523;
  wire wr_524;
  wire wr_525;
  wire wr_526;
  wire wr_527;
  wire wr_528;
  wire wr_529;
  wire wr_530;
  wire wr_531;
  wire wr_532;
  wire wr_533;
  wire wr_534;
  wire wr_535;
  wire wr_536;
  wire wr_537;
  wire wr_538;
  wire wr_539;
  wire wr_540;
  wire wr_541;
  wire wr_542;
  wire wr_543;
  wire wr_544;
  wire wr_545;
  wire wr_546;
  wire wr_547;
  wire wr_548;
  wire wr_549;
  wire wr_550;
  wire wr_551;
  wire wr_552;
  wire wr_553;
  wire wr_554;
  wire wr_555;
  wire wr_556;
  wire wr_557;
  wire wr_558;
  wire wr_559;
  wire wr_560;
  wire wr_561;
  wire wr_562;
  wire wr_563;
  wire wr_564;
  wire wr_565;
  wire wr_566;
  wire wr_567;
  wire wr_568;
  wire wr_569;
  wire wr_570;
  wire wr_571;
  wire wr_572;
  wire wr_573;
  wire wr_574;
  wire wr_575;
  wire wr_576;
  wire wr_577;
  wire wr_578;
  wire wr_579;
  wire wr_580;
  wire wr_581;
  wire wr_582;
  wire wr_583;
  wire wr_584;
  wire wr_585;
  wire wr_586;
  wire wr_587;
  wire wr_588;
  wire wr_589;
  wire wr_590;
  wire wr_591;
  wire wr_592;
  wire wr_593;
  wire wr_594;
  wire wr_595;
  wire wr_596;
  wire wr_597;
  wire wr_598;
  wire wr_599;
  wire wr_600;
  wire wr_601;
  wire wr_602;
  wire wr_603;
  wire wr_604;
  wire wr_605;
  wire wr_606;
  wire wr_607;
  wire wr_608;
  wire wr_609;
  wire wr_610;
  wire wr_611;
  wire wr_612;
  wire wr_613;
  wire wr_614;
  wire wr_615;
  wire wr_616;
  wire wr_617;
  wire wr_618;
  wire wr_619;
  wire wr_620;
  wire wr_621;
  wire wr_622;
  wire wr_623;
  wire wr_624;
  wire wr_625;
  wire wr_626;
  wire wr_627;
  wire wr_628;
  wire wr_629;
  wire wr_630;
  wire wr_631;
  wire wr_632;
  wire wr_633;
  wire wr_634;
  wire wr_635;
  wire wr_636;
  wire wr_637;
  wire wr_638;
  wire wr_639;
  wire wr_640;
  wire wr_641;
  wire wr_642;
  wire wr_643;
  wire wr_644;
  wire wr_645;
  wire wr_646;
  wire wr_647;
  wire wr_648;
  wire wr_649;
  wire wr_650;
  wire wr_651;
  wire wr_652;
  wire wr_653;
  wire wr_654;
  wire wr_655;
  wire wr_656;
  wire wr_657;
  wire wr_658;
  wire wr_659;
  wire wr_660;
  wire wr_661;
  wire wr_662;
  wire wr_663;
  wire wr_664;
  wire wr_665;
  wire wr_666;
  wire wr_667;
  wire wr_668;
  wire wr_669;
  wire wr_670;
  wire wr_671;
  wire wr_672;
  wire wr_673;
  wire wr_674;
  wire wr_675;
  wire wr_676;
  wire wr_677;
  wire wr_678;
  wire wr_679;
  wire wr_680;
  wire wr_681;
  wire wr_682;
  wire wr_683;
  wire wr_684;
  wire wr_685;
  wire wr_686;
  wire wr_687;
  wire wr_688;
  wire wr_689;
  wire wr_690;
  wire wr_691;
  wire wr_692;
  wire wr_693;
  wire wr_694;
  wire wr_695;
  wire wr_696;
  wire wr_697;
  wire wr_698;
  wire wr_699;
  wire wr_700;
  wire wr_701;
  wire wr_702;
  wire wr_703;
  wire wr_704;
  wire wr_705;
  wire wr_706;
  wire wr_707;
  wire wr_708;
  wire wr_709;
  wire wr_710;
  wire wr_711;
  wire wr_712;
  wire wr_713;
  wire wr_714;
  wire wr_715;
  wire wr_716;
  wire wr_717;
  wire wr_718;
  wire wr_719;
  wire wr_720;
  wire wr_721;
  wire wr_722;
  wire wr_723;
  wire wr_724;
  wire wr_725;
  wire wr_726;
  wire wr_727;
  wire wr_728;
  wire wr_729;
  wire wr_730;
  wire wr_731;
  wire wr_732;
  wire wr_733;
  wire wr_734;
  wire wr_735;
  wire wr_736;
  wire wr_737;
  wire wr_738;
  wire wr_739;
  wire wr_740;
  wire wr_741;
  wire wr_742;
  wire wr_743;
  wire wr_744;
  wire wr_745;
  wire wr_746;
  wire wr_747;
  wire wr_748;
  wire wr_749;
  wire wr_750;
  wire wr_751;
  wire wr_752;
  wire wr_753;
  wire wr_754;
  wire wr_755;
  wire wr_756;
  wire wr_757;
  wire wr_758;
  wire wr_759;
  wire wr_760;
  wire wr_761;
  wire wr_762;
  wire wr_763;
  wire wr_764;
  wire wr_765;
  wire wr_766;
  wire wr_767;
  wire wr_768;
  wire wr_769;
  wire wr_770;
  wire wr_771;
  wire wr_772;
  wire wr_773;
  wire wr_774;
  wire wr_775;
  wire wr_776;
  wire wr_777;
  wire wr_778;
  wire wr_779;
  wire wr_780;
  wire wr_781;
  wire wr_782;
  wire wr_783;
  wire wr_784;
  wire wr_785;
  wire wr_786;
  wire wr_787;
  wire wr_788;
  wire wr_789;
  wire wr_790;
  wire wr_791;
  wire wr_792;
  wire wr_793;
  wire wr_794;
  wire wr_795;
  wire wr_796;
  wire wr_797;
  wire wr_798;
  wire wr_799;
  wire wr_800;
  wire wr_801;
  wire wr_802;
  wire wr_803;
  wire wr_804;
  wire wr_805;
  wire wr_806;
  wire wr_807;
  wire wr_808;
  wire wr_809;
  wire wr_810;
  wire wr_811;
  wire wr_812;
  wire wr_813;
  wire wr_814;
  wire wr_815;
  wire wr_816;
  wire wr_817;
  wire wr_818;
  wire wr_819;
  wire wr_820;
  wire wr_821;
  wire wr_822;
  wire wr_823;
  wire wr_824;
  wire wr_825;
  wire wr_826;
  wire wr_827;
  wire wr_828;
  wire wr_829;
  wire wr_830;
  wire wr_831;
  wire wr_832;
  wire wr_833;
  wire wr_834;
  wire wr_835;
  wire wr_836;
  wire wr_837;
  wire wr_838;
  wire wr_839;
  wire wr_840;
  wire wr_841;
  wire wr_842;
  wire wr_843;
  wire wr_844;
  wire wr_845;
  wire wr_846;
  wire wr_847;
  wire wr_848;
  wire wr_849;
  wire wr_850;
  wire wr_851;
  wire wr_852;
  wire wr_853;
  wire wr_854;
  wire wr_855;
  wire wr_856;
  wire wr_857;
  wire wr_858;
  wire wr_859;
  wire wr_860;
  wire wr_861;
  wire wr_862;
  wire wr_863;
  wire wr_864;
  wire wr_865;
  wire wr_866;
  wire wr_867;
  wire wr_868;
  wire wr_869;
  wire wr_870;
  wire wr_871;
  wire wr_872;
  wire wr_873;
  wire wr_874;
  wire wr_875;
  wire wr_876;
  wire wr_877;
  wire wr_878;
  wire wr_879;
  wire wr_880;
  wire wr_881;
  wire wr_882;
  wire wr_883;
  wire wr_884;
  wire wr_885;
  wire wr_886;
  wire wr_887;
  wire wr_888;
  wire wr_889;
  wire wr_890;
  wire wr_891;
  wire wr_892;
  wire wr_893;
  wire wr_894;
  wire wr_895;
  wire wr_896;
  wire wr_897;
  wire wr_898;
  wire wr_899;
  wire wr_900;
  wire wr_901;
  wire wr_902;
  wire wr_903;
  wire wr_904;
  wire wr_905;
  wire wr_906;
  wire wr_907;
  wire wr_908;
  wire wr_909;
  wire wr_910;
  wire wr_911;
  wire wr_912;
  wire wr_913;
  wire wr_914;
  wire wr_915;
  wire wr_916;
  wire wr_917;
  wire wr_918;
  wire wr_919;
  wire wr_920;
  wire wr_921;
  wire wr_922;
  wire wr_923;
  wire wr_924;
  wire wr_925;
  wire wr_926;
  wire wr_927;
  wire wr_928;
  wire wr_929;
  wire wr_930;
  wire wr_931;
  wire wr_932;
  wire wr_933;
  wire wr_934;
  wire wr_935;
  wire wr_936;
  wire wr_937;
  wire wr_938;
  wire wr_939;
  wire wr_940;
  wire wr_941;
  wire wr_942;
  wire wr_943;
  wire wr_944;
  wire wr_945;
  wire wr_946;
  wire wr_947;
  wire wr_948;
  wire wr_949;
  wire wr_950;
  wire wr_951;
  wire wr_952;
  wire wr_953;
  wire wr_954;
  wire wr_955;
  wire wr_956;
  wire wr_957;
  wire wr_958;
  wire wr_959;
  wire wr_960;
  wire wr_961;
  wire wr_962;
  wire wr_963;
  wire wr_964;
  wire wr_965;
  wire wr_966;
  wire wr_967;
  wire wr_968;
  wire wr_969;
  wire wr_970;
  wire wr_971;
  wire wr_972;
  wire wr_973;
  wire wr_974;
  wire wr_975;
  wire wr_976;
  wire wr_977;
  wire wr_978;
  wire wr_979;
  wire wr_980;
  wire wr_981;
  wire wr_982;
  wire wr_983;
  wire wr_984;
  wire wr_985;
  wire wr_986;
  wire wr_987;
  wire wr_988;
  wire wr_989;
  wire wr_990;
  wire wr_991;
  wire wr_992;
  wire wr_993;
  wire wr_994;
  wire wr_995;
  wire wr_996;
  wire wr_997;
  wire wr_998;
  wire wr_999;
  wire wr_1000;
  wire wr_1001;
  wire wr_1002;
  wire wr_1003;
  wire wr_1004;
  wire wr_1005;
  wire wr_1006;
  wire wr_1007;
  wire wr_1008;
  wire wr_1009;
  wire wr_1010;
  wire wr_1011;
  wire wr_1012;
  wire wr_1013;
  wire wr_1014;
  wire wr_1015;
  wire wr_1016;
  wire wr_1017;
  wire wr_1018;
  wire wr_1019;
  wire wr_1020;
  wire wr_1021;
  wire wr_1022;
  wire wr_1023;
  wire wr_1024;
  wire wr_1025;
  wire wr_1026;
  wire wr_1027;
  wire wr_1028;
  wire wr_1029;
  wire wr_1030;
  wire wr_1031;
  wire wr_1032;
  wire wr_1033;
  wire wr_1034;
  wire wr_1035;
  wire wr_1036;
  wire wr_1037;
  wire wr_1038;
  wire wr_1039;
  wire wr_1040;
  wire wr_1041;
  wire wr_1042;
  wire wr_1043;
  wire wr_1044;
  wire wr_1045;
  wire wr_1046;
  wire wr_1047;
  wire wr_1048;
  wire wr_1049;
  wire wr_1050;
  wire wr_1051;
  wire wr_1052;
  wire wr_1053;
  wire wr_1054;
  wire wr_1055;
  wire wr_1056;
  wire wr_1057;
  wire wr_1058;
  wire wr_1059;
  wire wr_1060;
  wire wr_1061;
  wire wr_1062;
  wire wr_1063;
  wire wr_1064;
  wire wr_1065;
  wire wr_1066;
  wire wr_1067;
  wire wr_1068;
  wire wr_1069;
  wire wr_1070;
  wire wr_1071;
  wire wr_1072;
  wire wr_1073;
  wire wr_1074;
  wire wr_1075;
  wire wr_1076;
  wire wr_1077;
  wire wr_1078;
  wire wr_1079;
  wire wr_1080;
  wire wr_1081;
  wire wr_1082;
  wire wr_1083;
  wire wr_1084;
  wire wr_1085;
  wire wr_1086;
  wire wr_1087;
  wire wr_1088;
  wire wr_1089;
  wire wr_1090;
  wire wr_1091;
  wire wr_1092;
  wire wr_1093;
  wire wr_1094;
  wire wr_1095;
  wire wr_1096;
  wire wr_1097;
  wire wr_1098;
  wire wr_1099;
  wire wr_1100;
  wire wr_1101;
  wire wr_1102;
  wire wr_1103;
  wire wr_1104;
  wire wr_1105;
  wire wr_1106;
  wire wr_1107;
  wire wr_1108;
  wire wr_1109;
  wire wr_1110;
  wire wr_1111;
  wire wr_1112;
  wire wr_1113;
  wire wr_1114;
  wire wr_1115;
  wire wr_1116;
  wire wr_1117;
  wire wr_1118;
  wire wr_1119;
  wire wr_1120;
  wire wr_1121;
  wire wr_1122;
  wire wr_1123;
  wire wr_1124;
  wire wr_1125;
  wire wr_1126;
  wire wr_1127;
  wire wr_1128;
  wire wr_1129;
  wire wr_1130;
  wire wr_1131;
  wire wr_1132;
  wire wr_1133;
  wire wr_1134;
  wire wr_1135;
  wire wr_1136;
  wire wr_1137;
  wire wr_1138;
  wire wr_1139;
  wire wr_1140;
  wire wr_1141;
  wire wr_1142;
  wire wr_1143;
  wire wr_1144;
  wire wr_1145;
  wire wr_1146;
  wire wr_1147;
  wire wr_1148;
  wire wr_1149;
  wire wr_1150;
  wire wr_1151;
  wire wr_1152;
  wire wr_1153;
  wire wr_1154;
  wire wr_1155;
  wire wr_1156;
  wire wr_1157;
  wire wr_1158;
  wire wr_1159;
  wire wr_1160;
  wire wr_1161;
  wire wr_1162;
  wire wr_1163;
  wire wr_1164;
  wire wr_1165;
  wire wr_1166;
  wire wr_1167;
  wire wr_1168;
  wire wr_1169;
  wire wr_1170;
  wire wr_1171;
  wire wr_1172;
  wire wr_1173;
  wire wr_1174;
  wire wr_1175;
  wire wr_1176;
  wire wr_1177;
  wire wr_1178;
  wire wr_1179;
  wire wr_1180;
  wire wr_1181;
  wire wr_1182;
  wire wr_1183;
  wire wr_1184;
  wire wr_1185;
  wire wr_1186;
  wire wr_1187;
  wire wr_1188;
  wire wr_1189;
  wire wr_1190;
  wire wr_1191;
  wire wr_1192;
  wire wr_1193;
  wire wr_1194;
  wire wr_1195;
  wire wr_1196;
  wire wr_1197;
  wire wr_1198;
  wire wr_1199;
  wire wr_1200;
  wire wr_1201;
  wire wr_1202;
  wire wr_1203;
  wire wr_1204;
  wire wr_1205;
  wire wr_1206;
  wire wr_1207;
  wire wr_1208;
  wire wr_1209;
  wire wr_1210;
  wire wr_1211;
  wire wr_1212;
  wire wr_1213;
  wire wr_1214;
  wire wr_1215;
  wire wr_1216;
  wire wr_1217;
  wire wr_1218;
  wire wr_1219;
  wire wr_1220;
  wire wr_1221;
  wire wr_1222;
  wire wr_1223;
  wire wr_1224;
  wire wr_1225;
  wire wr_1226;
  wire wr_1227;
  wire wr_1228;
  wire wr_1229;
  wire wr_1230;
  wire wr_1231;
  wire wr_1232;
  wire wr_1233;
  wire wr_1234;
  wire wr_1235;
  wire wr_1236;
  wire wr_1237;
  wire wr_1238;
  wire wr_1239;
  wire wr_1240;
  wire wr_1241;
  wire wr_1242;
  wire wr_1243;
  wire wr_1244;
  wire wr_1245;
  wire wr_1246;
  wire wr_1247;
  wire wr_1248;
  wire wr_1249;
  wire wr_1250;
  wire wr_1251;
  wire wr_1252;
  wire wr_1253;
  wire wr_1254;
  wire wr_1255;
  wire wr_1256;
  wire wr_1257;
  wire wr_1258;
  wire wr_1259;
  wire wr_1260;
  wire wr_1261;
  wire wr_1262;
  wire wr_1263;
  wire wr_1264;
  wire wr_1265;
  wire wr_1266;
  wire wr_1267;
  wire wr_1268;
  wire wr_1269;
  wire wr_1270;
  wire wr_1271;
  wire wr_1272;
  wire wr_1273;
  wire wr_1274;
  wire wr_1275;
  wire wr_1276;
  wire wr_1277;
  wire wr_1278;
  wire wr_1279;
  wire wr_1280;
  wire wr_1281;
  wire wr_1282;
  wire wr_1283;
  wire wr_1284;
  wire wr_1285;
  wire wr_1286;
  wire wr_1287;
  wire wr_1288;
  wire wr_1289;
  wire wr_1290;
  wire wr_1291;
  wire wr_1292;
  wire wr_1293;
  wire wr_1294;
  wire wr_1295;
  wire wr_1296;
  wire wr_1297;
  wire wr_1298;
  wire wr_1299;
  wire wr_1300;
  wire wr_1301;
  wire wr_1302;
  wire wr_1303;
  wire wr_1304;
  wire wr_1305;
  wire wr_1306;
  wire wr_1307;
  wire wr_1308;
  wire wr_1309;
  wire wr_1310;
  wire wr_1311;
  wire wr_1312;
  wire wr_1313;
  wire wr_1314;
  wire wr_1315;
  wire wr_1316;
  wire wr_1317;
  wire wr_1318;
  wire wr_1319;
  wire wr_1320;
  wire wr_1321;
  wire wr_1322;
  wire wr_1323;
  wire wr_1324;
  wire wr_1325;
  wire wr_1326;
  wire wr_1327;
  wire wr_1328;
  wire wr_1329;
  wire wr_1330;
  wire wr_1331;
  wire wr_1332;
  wire wr_1333;
  wire wr_1334;
  wire wr_1335;
  wire wr_1336;
  wire wr_1337;
  wire wr_1338;
  wire wr_1339;
  wire wr_1340;
  wire wr_1341;
  wire wr_1342;
  wire wr_1343;
  wire wr_1344;
  wire wr_1345;
  wire wr_1346;
  wire wr_1347;
  wire wr_1348;
  wire wr_1349;
  wire wr_1350;
  wire wr_1351;
  wire wr_1352;
  wire wr_1353;
  wire wr_1354;
  wire wr_1355;
  wire wr_1356;
  wire wr_1357;
  wire wr_1358;
  wire wr_1359;
  wire wr_1360;
  wire wr_1361;
  wire wr_1362;
  wire wr_1363;
  wire wr_1364;
  wire wr_1365;
  wire wr_1366;
  wire wr_1367;
  wire wr_1368;
  wire wr_1369;
  wire wr_1370;
  wire wr_1371;
  wire wr_1372;
  wire wr_1373;
  wire wr_1374;
  wire wr_1375;
  wire wr_1376;
  wire wr_1377;
  wire wr_1378;
  wire wr_1379;
  wire wr_1380;
  wire wr_1381;
  wire wr_1382;
  wire wr_1383;
  wire wr_1384;
  wire wr_1385;
  wire wr_1386;
  wire wr_1387;
  wire wr_1388;
  wire wr_1389;
  wire wr_1390;
  wire wr_1391;
  wire wr_1392;
  wire wr_1393;
  wire wr_1394;
  wire wr_1395;
  wire wr_1396;
  wire wr_1397;
  wire wr_1398;
  wire wr_1399;
  wire wr_1400;
  wire wr_1401;
  wire wr_1402;
  wire wr_1403;
  wire wr_1404;
  wire wr_1405;
  wire wr_1406;
  wire wr_1407;
  wire wr_1408;
  wire wr_1409;
  wire wr_1410;
  wire wr_1411;
  wire wr_1412;
  wire wr_1413;
  wire wr_1414;
  wire wr_1415;
  wire wr_1416;
  wire wr_1417;
  wire wr_1418;
  wire wr_1419;
  wire wr_1420;
  wire wr_1421;
  wire wr_1422;
  wire wr_1423;
  wire wr_1424;
  wire wr_1425;
  wire wr_1426;
  wire wr_1427;
  wire wr_1428;
  wire wr_1429;
  wire wr_1430;
  wire wr_1431;
  wire wr_1432;
  wire wr_1433;
  wire wr_1434;
  wire wr_1435;
  wire wr_1436;
  wire wr_1437;
  wire wr_1438;
  wire wr_1439;
  wire wr_1440;
  wire wr_1441;
  wire wr_1442;
  wire wr_1443;
  wire wr_1444;
  wire wr_1445;
  wire wr_1446;
  wire wr_1447;
  wire wr_1448;
  wire wr_1449;
  wire wr_1450;
  wire wr_1451;
  wire wr_1452;
  wire wr_1453;
  wire wr_1454;
  wire wr_1455;
  wire wr_1456;
  wire wr_1457;
  wire wr_1458;
  wire wr_1459;
  wire wr_1460;
  wire wr_1461;
  wire wr_1462;
  wire wr_1463;
  wire wr_1464;
  wire wr_1465;
  wire wr_1466;
  wire wr_1467;
  wire wr_1468;
  wire wr_1469;
  wire wr_1470;
  wire wr_1471;
  wire wr_1472;
  wire wr_1473;
  wire wr_1474;
  wire wr_1475;
  wire wr_1476;
  wire wr_1477;
  wire wr_1478;
  wire wr_1479;
  wire wr_1480;
  wire wr_1481;
  wire wr_1482;
  wire wr_1483;
  wire wr_1484;
  wire wr_1485;
  wire wr_1486;
  wire wr_1487;
  wire wr_1488;
  wire wr_1489;
  wire wr_1490;
  wire wr_1491;
  wire wr_1492;
  wire wr_1493;
  wire wr_1494;
  wire wr_1495;
  wire wr_1496;
  wire wr_1497;
  wire wr_1498;
  wire wr_1499;
  wire wr_1500;
  wire wr_1501;
  wire wr_1502;
  wire wr_1503;
  wire wr_1504;
  wire wr_1505;
  wire wr_1506;
  wire wr_1507;
  wire wr_1508;
  wire wr_1509;
  wire wr_1510;
  wire wr_1511;
  wire wr_1512;
  wire wr_1513;
  wire wr_1514;
  wire wr_1515;
  wire wr_1516;
  wire wr_1517;
  wire wr_1518;
  wire wr_1519;
  wire wr_1520;
  wire wr_1521;
  wire wr_1522;
  wire wr_1523;
  wire wr_1524;
  wire wr_1525;
  wire wr_1526;
  wire wr_1527;
  wire wr_1528;
  wire wr_1529;
  wire wr_1530;
  wire wr_1531;
  wire wr_1532;
  wire wr_1533;
  wire wr_1534;
  wire wr_1535;
  wire wr_1536;
  wire wr_1537;
  wire wr_1538;
  wire wr_1539;
  wire wr_1540;
  wire wr_1541;
  wire wr_1542;
  wire wr_1543;
  wire wr_1544;
  wire wr_1545;
  wire wr_1546;
  wire wr_1547;
  wire wr_1548;
  wire wr_1549;
  wire wr_1550;
  wire wr_1551;
  wire wr_1552;
  wire wr_1553;
  wire wr_1554;
  wire wr_1555;
  wire wr_1556;
  wire wr_1557;
  wire wr_1558;
  wire wr_1559;
  wire wr_1560;
  wire wr_1561;
  wire wr_1562;
  wire wr_1563;
  wire wr_1564;
  wire wr_1565;
  wire wr_1566;
  wire wr_1567;
  wire wr_1568;
  wire wr_1569;
  wire wr_1570;
  wire wr_1571;
  wire wr_1572;
  wire wr_1573;
  wire wr_1574;
  wire wr_1575;
  wire wr_1576;
  wire wr_1577;
  wire wr_1578;
  wire wr_1579;
  wire wr_1580;
  wire wr_1581;
  wire wr_1582;
  wire wr_1583;
  wire wr_1584;
  wire wr_1585;
  wire wr_1586;
  wire wr_1587;
  wire wr_1588;
  wire wr_1589;
  wire wr_1590;
  wire wr_1591;
  wire wr_1592;
  wire wr_1593;
  wire wr_1594;
  wire wr_1595;
  wire wr_1596;
  wire wr_1597;
  wire wr_1598;
  wire wr_1599;
  wire wr_1600;
  wire wr_1601;
  wire wr_1602;
  wire wr_1603;
  wire wr_1604;
  wire wr_1605;
  wire wr_1606;
  wire wr_1607;
  wire wr_1608;
  wire wr_1609;
  wire wr_1610;
  wire wr_1611;
  wire wr_1612;
  wire wr_1613;
  wire wr_1614;
  wire wr_1615;
  wire wr_1616;
  wire wr_1617;
  wire wr_1618;
  wire wr_1619;
  wire wr_1620;
  wire wr_1621;
  wire wr_1622;
  wire wr_1623;
  wire wr_1624;
  wire wr_1625;
  wire wr_1626;
  wire wr_1627;
  wire wr_1628;
  wire wr_1629;
  wire wr_1630;
  wire wr_1631;
  wire wr_1632;
  wire wr_1633;
  wire wr_1634;
  wire wr_1635;
  wire wr_1636;
  wire wr_1637;
  wire wr_1638;
  wire wr_1639;
  wire wr_1640;
  wire wr_1641;
  wire wr_1642;
  wire wr_1643;
  wire wr_1644;
  wire wr_1645;
  wire wr_1646;
  wire wr_1647;
  wire wr_1648;
  wire wr_1649;
  wire wr_1650;
  wire wr_1651;
  wire wr_1652;
  wire wr_1653;
  wire wr_1654;
  wire wr_1655;
  wire wr_1656;
  wire wr_1657;
  wire wr_1658;
  wire wr_1659;
  wire wr_1660;
  wire wr_1661;
  wire wr_1662;
  wire wr_1663;
  wire wr_1664;
  wire wr_1665;
  wire wr_1666;
  wire wr_1667;
  wire wr_1668;
  wire wr_1669;
  wire wr_1670;
  wire wr_1671;
  wire wr_1672;
  wire wr_1673;
  wire wr_1674;
  wire wr_1675;
  wire wr_1676;
  wire wr_1677;
  wire wr_1678;
  wire wr_1679;
  wire wr_1680;
  wire wr_1681;
  wire wr_1682;
  wire wr_1683;
  wire wr_1684;
  wire wr_1685;
  wire wr_1686;
  wire wr_1687;
  wire wr_1688;
  wire wr_1689;
  wire wr_1690;
  wire wr_1691;
  wire wr_1692;
  wire wr_1693;
  wire wr_1694;
  wire wr_1695;
  wire wr_1696;
  wire wr_1697;
  wire wr_1698;
  wire wr_1699;
  wire wr_1700;
  wire wr_1701;
  wire wr_1702;
  wire wr_1703;
  wire wr_1704;
  wire wr_1705;
  wire wr_1706;
  wire wr_1707;
  wire wr_1708;
  wire wr_1709;
  wire wr_1710;
  wire wr_1711;
  wire wr_1712;
  wire wr_1713;
  wire wr_1714;
  wire wr_1715;
  wire wr_1716;
  wire wr_1717;
  wire wr_1718;
  wire wr_1719;
  wire wr_1720;
  wire wr_1721;
  wire wr_1722;
  wire wr_1723;
  wire wr_1724;
  wire wr_1725;
  wire wr_1726;
  wire wr_1727;
  wire wr_1728;
  wire wr_1729;
  wire wr_1730;
  wire wr_1731;
  wire wr_1732;
  wire wr_1733;
  wire wr_1734;
  wire wr_1735;
  wire wr_1736;
  wire wr_1737;
  wire wr_1738;
  wire wr_1739;
  wire wr_1740;
  wire wr_1741;
  wire wr_1742;
  wire wr_1743;
  wire wr_1744;
  wire wr_1745;
  wire wr_1746;
  wire wr_1747;
  wire wr_1748;
  wire wr_1749;
  wire wr_1750;
  wire wr_1751;
  wire wr_1752;
  wire wr_1753;
  wire wr_1754;
  wire wr_1755;
  wire wr_1756;
  wire wr_1757;
  wire wr_1758;
  wire wr_1759;
  wire wr_1760;
  wire wr_1761;
  wire wr_1762;
  wire wr_1763;
  wire wr_1764;
  wire wr_1765;
  wire wr_1766;
  wire wr_1767;
  wire wr_1768;
  wire wr_1769;
  wire wr_1770;
  wire wr_1771;
  wire wr_1772;
  wire wr_1773;
  wire wr_1774;
  wire wr_1775;
  wire wr_1776;
  wire wr_1777;
  wire wr_1778;
  wire wr_1779;
  wire wr_1780;
  wire wr_1781;
  wire wr_1782;
  wire wr_1783;
  wire wr_1784;
  wire wr_1785;
  wire wr_1786;
  wire wr_1787;
  wire wr_1788;
  wire wr_1789;
  wire wr_1790;
  wire wr_1791;
  wire wr_1792;
  wire wr_1793;
  wire wr_1794;
  wire wr_1795;
  wire wr_1796;
  wire wr_1797;
  wire wr_1798;
  wire wr_1799;
  wire wr_1800;
  wire wr_1801;
  wire wr_1802;
  wire wr_1803;
  wire wr_1804;
  wire wr_1805;
  wire wr_1806;
  wire wr_1807;
  wire wr_1808;
  wire wr_1809;
  wire wr_1810;
  wire wr_1811;
  wire wr_1812;
  wire wr_1813;
  wire wr_1814;
  wire wr_1815;
  wire wr_1816;
  wire wr_1817;
  wire wr_1818;
  wire wr_1819;
  wire wr_1820;
  wire wr_1821;
  wire wr_1822;
  wire wr_1823;
  wire wr_1824;
  wire wr_1825;
  wire wr_1826;
  wire wr_1827;
  wire wr_1828;
  wire wr_1829;
  wire wr_1830;
  wire wr_1831;
  wire wr_1832;
  wire wr_1833;
  wire wr_1834;
  wire wr_1835;
  wire wr_1836;
  wire wr_1837;
  wire wr_1838;
  wire wr_1839;
  wire wr_1840;
  wire wr_1841;
  wire wr_1842;
  wire wr_1843;
  wire wr_1844;
  wire wr_1845;
  wire wr_1846;
  wire wr_1847;
  wire wr_1848;
  wire wr_1849;
  wire wr_1850;
  wire wr_1851;
  wire wr_1852;
  wire wr_1853;
  wire wr_1854;
  wire wr_1855;
  wire wr_1856;
  wire wr_1857;
  wire wr_1858;
  wire wr_1859;
  wire wr_1860;
  wire wr_1861;
  wire wr_1862;
  wire wr_1863;
  wire wr_1864;
  wire wr_1865;
  wire wr_1866;
  wire wr_1867;
  wire wr_1868;
  wire wr_1869;
  wire wr_1870;
  wire wr_1871;
  wire wr_1872;
  wire wr_1873;
  wire wr_1874;
  wire wr_1875;
  wire wr_1876;
  wire wr_1877;
  wire wr_1878;
  wire wr_1879;
  wire wr_1880;
  wire wr_1881;
  wire wr_1882;
  wire wr_1883;
  wire wr_1884;
  wire wr_1885;
  wire wr_1886;
  wire wr_1887;
  wire wr_1888;
  wire wr_1889;
  wire wr_1890;
  wire wr_1891;
  wire wr_1892;
  wire wr_1893;
  wire wr_1894;
  wire wr_1895;
  wire wr_1896;
  wire wr_1897;
  wire wr_1898;
  wire wr_1899;
  wire wr_1900;
  wire wr_1901;
  wire wr_1902;
  wire wr_1903;
  wire wr_1904;
  wire wr_1905;
  wire wr_1906;
  wire wr_1907;
  wire wr_1908;
  wire wr_1909;
  wire wr_1910;
  wire wr_1911;
  wire wr_1912;
  wire wr_1913;
  wire wr_1914;
  wire wr_1915;
  wire wr_1916;
  wire wr_1917;
  wire wr_1918;
  wire wr_1919;
  wire wr_1920;
  wire wr_1921;
  wire wr_1922;
  wire wr_1923;
  wire wr_1924;
  wire wr_1925;
  wire wr_1926;
  wire wr_1927;
  wire wr_1928;
  wire wr_1929;
  wire wr_1930;
  wire wr_1931;
  wire wr_1932;
  wire wr_1933;
  wire wr_1934;
  wire wr_1935;
  wire wr_1936;
  wire wr_1937;
  wire wr_1938;
  wire wr_1939;
  wire wr_1940;
  wire wr_1941;
  wire wr_1942;
  wire wr_1943;
  wire wr_1944;
  wire wr_1945;
  wire wr_1946;
  wire wr_1947;
  wire wr_1948;
  wire wr_1949;
  wire wr_1950;
  wire wr_1951;
  wire wr_1952;
  wire wr_1953;
  wire wr_1954;
  wire wr_1955;
  wire wr_1956;
  wire wr_1957;
  wire wr_1958;
  wire wr_1959;
  wire wr_1960;
  wire wr_1961;
  wire wr_1962;
  wire wr_1963;
  wire wr_1964;
  wire wr_1965;
  wire wr_1966;
  wire wr_1967;
  wire wr_1968;
  wire wr_1969;
  wire wr_1970;
  wire wr_1971;
  wire wr_1972;
  wire wr_1973;
  wire wr_1974;
  wire wr_1975;
  wire wr_1976;
  wire wr_1977;
  wire wr_1978;
  wire wr_1979;
  wire wr_1980;
  wire wr_1981;
  wire wr_1982;
  wire wr_1983;
  wire wr_1984;
  wire wr_1985;
  wire wr_1986;
  wire wr_1987;
  wire wr_1988;
  wire wr_1989;
  wire wr_1990;
  wire wr_1991;
  wire wr_1992;
  wire wr_1993;
  wire wr_1994;
  wire wr_1995;
  wire wr_1996;
  wire wr_1997;
  wire wr_1998;
  wire wr_1999;
  wire wr_2000;
  wire wr_2001;
  wire wr_2002;
  wire wr_2003;
  wire wr_2004;
  wire wr_2005;
  wire wr_2006;
  wire wr_2007;
  wire wr_2008;
  wire wr_2009;
  wire wr_2010;
  wire wr_2011;
  wire wr_2012;
  wire wr_2013;
  wire wr_2014;
  wire wr_2015;
  wire wr_2016;
  wire wr_2017;
  wire wr_2018;
  wire wr_2019;
  wire wr_2020;
  wire wr_2021;
  wire wr_2022;
  wire wr_2023;
  wire wr_2024;
  wire wr_2025;
  wire wr_2026;
  wire wr_2027;
  wire wr_2028;
  wire wr_2029;
  wire wr_2030;
  wire wr_2031;
  wire wr_2032;
  wire wr_2033;
  wire wr_2034;
  wire wr_2035;
  wire wr_2036;
  wire wr_2037;
  wire wr_2038;
  wire wr_2039;
  wire wr_2040;
  wire wr_2041;
  wire wr_2042;
  wire wr_2043;
  wire wr_2044;
  wire wr_2045;
  wire wr_2046;
  wire wr_2047;
  wire wr_2048;
  wire wr_2049;
  wire wr_2050;
  wire wr_2051;
  wire wr_2052;
  wire wr_2053;
  wire wr_2054;
  wire wr_2055;
  wire wr_2056;
  wire wr_2057;
  wire wr_2058;
  wire wr_2059;
  wire wr_2060;
  wire wr_2061;
  wire wr_2062;
  wire wr_2063;
  wire wr_2064;
  wire wr_2065;
  wire wr_2066;
  wire wr_2067;
  wire wr_2068;
  wire wr_2069;
  wire wr_2070;
  wire wr_2071;
  wire wr_2072;
  wire wr_2073;
  wire wr_2074;
  wire wr_2075;
  wire wr_2076;
  wire wr_2077;
  wire wr_2078;
  wire wr_2079;
  wire wr_2080;
  wire wr_2081;
  wire wr_2082;
  wire wr_2083;
  wire wr_2084;
  wire wr_2085;
  wire wr_2086;
  wire wr_2087;
  wire wr_2088;
  wire wr_2089;
  wire wr_2090;
  wire wr_2091;
  wire wr_2092;
  wire wr_2093;
  wire wr_2094;
  wire wr_2095;
  wire wr_2096;
  wire wr_2097;
  wire wr_2098;
  wire wr_2099;
  wire wr_2100;
  wire wr_2101;
  wire wr_2102;
  wire wr_2103;
  wire wr_2104;
  wire wr_2105;
  wire wr_2106;
  wire wr_2107;
  wire wr_2108;
  wire wr_2109;
  wire wr_2110;
  wire wr_2111;
  wire wr_2112;
  wire wr_2113;
  wire wr_2114;
  wire wr_2115;
  wire wr_2116;
  wire wr_2117;
  wire wr_2118;
  wire wr_2119;
  wire wr_2120;
  wire wr_2121;
  wire wr_2122;
  wire wr_2123;
  wire wr_2124;
  wire wr_2125;
  wire wr_2126;
  wire wr_2127;
  wire wr_2128;
  wire wr_2129;
  wire wr_2130;
  wire wr_2131;
  wire wr_2132;
  wire wr_2133;
  wire wr_2134;
  wire wr_2135;
  wire wr_2136;
  wire wr_2137;
  wire wr_2138;
  wire wr_2139;
  wire wr_2140;
  wire wr_2141;
  wire wr_2142;
  wire wr_2143;
  wire wr_2144;
  wire wr_2145;
  wire wr_2146;
  wire wr_2147;
  wire wr_2148;
  wire wr_2149;
  wire wr_2150;
  wire wr_2151;
  wire wr_2152;
  wire wr_2153;
  wire wr_2154;
  wire wr_2155;
  wire wr_2156;
  wire wr_2157;
  wire wr_2158;
  wire wr_2159;
  wire wr_2160;
  wire wr_2161;
  wire wr_2162;
  wire wr_2163;
  wire wr_2164;
  wire wr_2165;
  wire wr_2166;
  wire wr_2167;
  wire wr_2168;
  wire wr_2169;
  wire wr_2170;
  wire wr_2171;
  wire wr_2172;
  wire wr_2173;
  wire wr_2174;
  wire wr_2175;
  wire wr_2176;
  wire wr_2177;
  wire wr_2178;
  wire wr_2179;
  wire wr_2180;
  wire wr_2181;
  wire wr_2182;
  wire wr_2183;
  wire wr_2184;
  wire wr_2185;
  wire wr_2186;
  wire wr_2187;
  wire wr_2188;
  wire wr_2189;
  wire wr_2190;
  wire wr_2191;
  wire wr_2192;
  wire wr_2193;
  wire wr_2194;
  wire wr_2195;
  wire wr_2196;
  wire wr_2197;
  wire wr_2198;
  wire wr_2199;
  wire wr_2200;
  wire wr_2201;
  wire wr_2202;
  wire wr_2203;
  wire wr_2204;
  wire wr_2205;
  wire wr_2206;
  wire wr_2207;
  wire wr_2208;
  wire wr_2209;
  wire wr_2210;
  wire wr_2211;
  wire wr_2212;
  wire wr_2213;
  wire wr_2214;
  wire wr_2215;
  wire wr_2216;
  wire wr_2217;
  wire wr_2218;
  wire wr_2219;
  wire wr_2220;
  wire wr_2221;
  wire wr_2222;
  wire wr_2223;
  wire wr_2224;
  wire wr_2225;
  wire wr_2226;
  wire wr_2227;
  wire wr_2228;
  wire wr_2229;
  wire wr_2230;
  wire wr_2231;
  wire wr_2232;
  wire wr_2233;
  wire wr_2234;
  wire wr_2235;
  wire wr_2236;
  wire wr_2237;
  wire wr_2238;
  wire wr_2239;
  wire wr_2240;
  wire wr_2241;
  wire wr_2242;
  wire wr_2243;
  wire wr_2244;
  wire wr_2245;
  wire wr_2246;
  wire wr_2247;
  wire wr_2248;
  wire wr_2249;
  wire wr_2250;
  wire wr_2251;
  wire wr_2252;
  wire wr_2253;
  wire wr_2254;
  wire wr_2255;
  wire wr_2256;
  wire wr_2257;
  wire wr_2258;
  wire wr_2259;
  wire wr_2260;
  wire wr_2261;
  wire wr_2262;
  wire wr_2263;
  wire wr_2264;
  wire wr_2265;
  wire wr_2266;
  wire wr_2267;
  wire wr_2268;
  wire wr_2269;
  wire wr_2270;
  wire wr_2271;
  wire wr_2272;
  wire wr_2273;
  wire wr_2274;
  wire wr_2275;
  wire wr_2276;
  wire wr_2277;
  wire wr_2278;
  wire wr_2279;
  wire wr_2280;
  wire wr_2281;
  wire wr_2282;
  wire wr_2283;
  wire wr_2284;
  wire wr_2285;
  wire wr_2286;
  wire wr_2287;
  wire wr_2288;
  wire wr_2289;
  wire wr_2290;
  wire wr_2291;
  wire wr_2292;
  wire wr_2293;
  wire wr_2294;
  wire wr_2295;
  wire wr_2296;
  wire wr_2297;
  wire wr_2298;
  wire wr_2299;
  wire wr_2300;
  wire wr_2301;
  wire wr_2302;
  wire wr_2303;
  wire wr_2304;
  wire wr_2305;
  wire wr_2306;
  wire wr_2307;
  wire wr_2308;
  wire wr_2309;
  wire wr_2310;
  wire wr_2311;
  wire wr_2312;
  wire wr_2313;
  wire wr_2314;
  wire wr_2315;
  wire wr_2316;
  wire wr_2317;
  wire wr_2318;
  wire wr_2319;
  wire wr_2320;
  wire wr_2321;
  wire wr_2322;
  wire wr_2323;
  wire wr_2324;
  wire wr_2325;
  wire wr_2326;
  wire wr_2327;
  wire wr_2328;
  wire wr_2329;
  wire wr_2330;
  wire wr_2331;
  wire wr_2332;
  wire wr_2333;
  wire wr_2334;
  wire wr_2335;
  wire wr_2336;
  wire wr_2337;
  wire wr_2338;
  wire wr_2339;
  wire wr_2340;
  wire wr_2341;
  wire wr_2342;
  wire wr_2343;
  wire wr_2344;
  wire wr_2345;
  wire wr_2346;
  wire wr_2347;
  wire wr_2348;
  wire wr_2349;
  wire wr_2350;
  wire wr_2351;
  wire wr_2352;
  wire wr_2353;
  wire wr_2354;
  wire wr_2355;
  wire wr_2356;
  wire wr_2357;
  wire wr_2358;
  wire wr_2359;
  wire wr_2360;
  wire wr_2361;
  wire wr_2362;
  wire wr_2363;
  wire wr_2364;
  wire wr_2365;
  wire wr_2366;
  wire wr_2367;
  wire wr_2368;
  wire wr_2369;
  wire wr_2370;
  wire wr_2371;
  wire wr_2372;
  wire wr_2373;
  wire wr_2374;
  wire wr_2375;
  wire wr_2376;
  wire wr_2377;
  wire wr_2378;
  wire wr_2379;
  wire wr_2380;
  wire wr_2381;
  wire wr_2382;
  wire wr_2383;
  wire wr_2384;
  wire wr_2385;
  wire wr_2386;
  wire wr_2387;
  wire wr_2388;
  wire wr_2389;
  wire wr_2390;
  wire wr_2391;
  wire wr_2392;
  wire wr_2393;
  wire wr_2394;
  wire wr_2395;
  wire wr_2396;
  wire wr_2397;
  wire wr_2398;
  wire wr_2399;
  wire wr_2400;
  wire wr_2401;
  wire wr_2402;
  wire wr_2403;
  wire wr_2404;
  wire wr_2405;
  wire wr_2406;
  wire wr_2407;
  wire wr_2408;
  wire wr_2409;
  wire wr_2410;
  wire wr_2411;
  wire wr_2412;
  wire wr_2413;
  wire wr_2414;
  wire wr_2415;
  wire wr_2416;
  wire wr_2417;
  wire wr_2418;
  wire wr_2419;
  wire wr_2420;
  wire wr_2421;
  wire wr_2422;
  wire wr_2423;
  wire wr_2424;
  wire wr_2425;
  wire wr_2426;
  wire wr_2427;
  wire wr_2428;
  wire wr_2429;
  wire wr_2430;
  wire wr_2431;
  wire wr_2432;
  wire wr_2433;
  wire wr_2434;
  wire wr_2435;
  wire wr_2436;
  wire wr_2437;
  wire wr_2438;
  wire wr_2439;
  wire wr_2440;
  wire wr_2441;
  wire wr_2442;
  wire wr_2443;
  wire wr_2444;
  wire wr_2445;
  wire wr_2446;
  wire wr_2447;
  wire wr_2448;
  wire wr_2449;
  wire wr_2450;
  wire wr_2451;
  wire wr_2452;
  wire wr_2453;
  wire wr_2454;
  wire wr_2455;
  wire wr_2456;
  wire wr_2457;
  wire wr_2458;
  wire wr_2459;
  wire wr_2460;
  wire wr_2461;
  wire wr_2462;
  wire wr_2463;
  wire wr_2464;
  wire wr_2465;
  wire wr_2466;
  wire wr_2467;
  wire wr_2468;
  wire wr_2469;
  wire wr_2470;
  wire wr_2471;
  wire wr_2472;
  wire wr_2473;
  wire wr_2474;
  wire wr_2475;
  wire wr_2476;
  wire wr_2477;
  wire wr_2478;
  wire wr_2479;
  wire wr_2480;
  wire wr_2481;
  wire wr_2482;
  wire wr_2483;
  wire wr_2484;
  wire wr_2485;
  wire wr_2486;
  wire wr_2487;
  wire wr_2488;
  wire wr_2489;
  wire wr_2490;
  wire wr_2491;
  wire wr_2492;
  wire wr_2493;
  wire wr_2494;
  wire wr_2495;
  wire wr_2496;
  wire wr_2497;
  wire wr_2498;
  wire wr_2499;
  wire wr_2500;
  wire wr_2501;
  wire wr_2502;
  wire wr_2503;
  wire wr_2504;
  wire wr_2505;
  wire wr_2506;
  wire wr_2507;
  wire wr_2508;
  wire wr_2509;
  wire wr_2510;
  wire wr_2511;
  wire wr_2512;
  wire wr_2513;
  wire wr_2514;
  wire wr_2515;
  wire wr_2516;
  wire wr_2517;
  wire wr_2518;
  wire wr_2519;
  wire wr_2520;
  wire wr_2521;
  wire wr_2522;
  wire wr_2523;
  wire wr_2524;
  wire wr_2525;
  wire wr_2526;
  wire wr_2527;
  wire wr_2528;
  wire wr_2529;
  wire wr_2530;
  wire wr_2531;
  wire wr_2532;
  wire wr_2533;
  wire wr_2534;
  wire wr_2535;
  wire wr_2536;
  wire wr_2537;
  wire wr_2538;
  wire wr_2539;
  wire wr_2540;
  wire wr_2541;
  wire wr_2542;
  wire wr_2543;
  wire wr_2544;
  wire wr_2545;
  wire wr_2546;
  wire wr_2547;
  wire wr_2548;
  wire wr_2549;
  wire wr_2550;
  wire wr_2551;
  wire wr_2552;
  wire wr_2553;
  wire wr_2554;
  wire wr_2555;
  wire wr_2556;
  wire wr_2557;
  wire wr_2558;
  wire wr_2559;
  wire wr_2560;
  wire wr_2561;
  wire wr_2562;
  wire wr_2563;
  wire wr_2564;
  wire wr_2565;
  wire wr_2566;
  wire wr_2567;
  wire wr_2568;
  wire wr_2569;
  wire wr_2570;
  wire wr_2571;
  wire wr_2572;
  wire wr_2573;
  wire wr_2574;
  wire wr_2575;
  wire wr_2576;
  wire wr_2577;
  wire wr_2578;
  wire wr_2579;
  wire wr_2580;
  wire wr_2581;
  wire wr_2582;
  wire wr_2583;
  wire wr_2584;
  wire wr_2585;
  wire wr_2586;
  wire wr_2587;
  wire wr_2588;
  wire wr_2589;
  wire wr_2590;
  wire wr_2591;
  wire wr_2592;
  wire wr_2593;
  wire wr_2594;
  wire wr_2595;
  wire wr_2596;
  wire wr_2597;
  wire wr_2598;
  wire wr_2599;
  wire wr_2600;
  wire wr_2601;
  wire wr_2602;
  wire wr_2603;
  wire wr_2604;
  wire wr_2605;
  wire wr_2606;
  wire wr_2607;
  wire wr_2608;
  wire wr_2609;
  wire wr_2610;
  wire wr_2611;
  wire wr_2612;
  wire wr_2613;
  wire wr_2614;
  wire wr_2615;
  wire wr_2616;
  wire wr_2617;
  wire wr_2618;
  wire wr_2619;
  wire wr_2620;
  wire wr_2621;
  wire wr_2622;
  wire wr_2623;
  wire wr_2624;
  wire wr_2625;
  wire wr_2626;
  wire wr_2627;
  wire wr_2628;
  wire wr_2629;
  wire wr_2630;
  wire wr_2631;
  wire wr_2632;
  wire wr_2633;
  wire wr_2634;
  wire wr_2635;
  wire wr_2636;
  wire wr_2637;
  wire wr_2638;
  wire wr_2639;
  wire wr_2640;
  wire wr_2641;
  wire wr_2642;
  wire wr_2643;
  wire wr_2644;
  wire wr_2645;
  wire wr_2646;
  wire wr_2647;
  wire wr_2648;
  wire wr_2649;
  wire wr_2650;
  wire wr_2651;
  wire wr_2652;
  wire wr_2653;
  wire wr_2654;
  wire wr_2655;
  wire wr_2656;
  wire wr_2657;
  wire wr_2658;
  wire wr_2659;
  wire wr_2660;
  wire wr_2661;
  wire wr_2662;
  wire wr_2663;
  wire wr_2664;
  wire wr_2665;
  wire wr_2666;
  wire wr_2667;
  wire wr_2668;
  wire wr_2669;
  wire wr_2670;
  wire wr_2671;
  wire wr_2672;
  wire wr_2673;
  wire wr_2674;
  wire wr_2675;
  wire wr_2676;
  wire wr_2677;
  wire wr_2678;
  wire wr_2679;
  wire wr_2680;
  wire wr_2681;
  wire wr_2682;
  wire wr_2683;
  wire wr_2684;
  wire wr_2685;
  wire wr_2686;
  wire wr_2687;
  wire wr_2688;
  wire wr_2689;
  wire wr_2690;
  wire wr_2691;
  wire wr_2692;
  wire wr_2693;
  wire wr_2694;
  wire wr_2695;
  wire wr_2696;
  wire wr_2697;
  wire wr_2698;
  wire wr_2699;
  wire wr_2700;
  wire wr_2701;
  wire wr_2702;
  wire wr_2703;
  wire wr_2704;
  wire wr_2705;
  wire wr_2706;
  wire wr_2707;
  wire wr_2708;
  wire wr_2709;
  wire wr_2710;
  wire wr_2711;
  wire wr_2712;
  wire wr_2713;
  wire wr_2714;
  wire wr_2715;
  wire wr_2716;
  wire wr_2717;
  wire wr_2718;
  wire wr_2719;
  wire wr_2720;
  wire wr_2721;
  wire wr_2722;
  wire wr_2723;
  wire wr_2724;
  wire wr_2725;
  wire wr_2726;
  wire wr_2727;
  wire wr_2728;
  wire wr_2729;
  wire wr_2730;
  wire wr_2731;
  wire wr_2732;
  wire wr_2733;
  wire wr_2734;
  wire wr_2735;
  wire wr_2736;
  wire wr_2737;
  wire wr_2738;
  wire wr_2739;
  wire wr_2740;
  wire wr_2741;
  wire wr_2742;
  wire wr_2743;
  wire wr_2744;
  wire wr_2745;
  wire wr_2746;
  wire wr_2747;
  wire wr_2748;
  wire wr_2749;
  wire wr_2750;
  wire wr_2751;
  wire wr_2752;
  wire wr_2753;
  wire wr_2754;
  wire wr_2755;
  wire wr_2756;
  wire wr_2757;
  wire wr_2758;
  wire wr_2759;
  wire wr_2760;
  wire wr_2761;
  wire wr_2762;
  wire wr_2763;
  wire wr_2764;
  wire wr_2765;
  wire wr_2766;
  wire wr_2767;
  wire wr_2768;
  wire wr_2769;
  wire wr_2770;
  wire wr_2771;
  wire wr_2772;
  wire wr_2773;
  wire wr_2774;
  wire wr_2775;
  wire wr_2776;
  wire wr_2777;
  wire wr_2778;
  wire wr_2779;
  wire wr_2780;
  wire wr_2781;
  wire wr_2782;
  wire wr_2783;
  wire wr_2784;
  wire wr_2785;
  wire wr_2786;
  wire wr_2787;
  wire wr_2788;
  wire wr_2789;
  wire wr_2790;
  wire wr_2791;
  wire wr_2792;
  wire wr_2793;
  wire wr_2794;
  wire wr_2795;
  wire wr_2796;
  wire wr_2797;
  wire wr_2798;
  wire wr_2799;
  wire wr_2800;
  wire wr_2801;
  wire wr_2802;
  wire wr_2803;
  wire wr_2804;
  wire wr_2805;
  wire wr_2806;
  wire wr_2807;
  wire wr_2808;
  wire wr_2809;
  wire wr_2810;
  wire wr_2811;
  wire wr_2812;
  wire wr_2813;
  wire wr_2814;
  wire wr_2815;
  wire wr_2816;
  wire wr_2817;
  wire wr_2818;
  wire wr_2819;
  wire wr_2820;
  wire wr_2821;
  wire wr_2822;
  wire wr_2823;
  wire wr_2824;
  wire wr_2825;
  wire wr_2826;
  wire wr_2827;
  wire wr_2828;
  wire wr_2829;
  wire wr_2830;
  wire wr_2831;
  wire wr_2832;
  wire wr_2833;
  wire wr_2834;
  wire wr_2835;
  wire wr_2836;
  wire wr_2837;
  wire wr_2838;
  wire wr_2839;
  wire wr_2840;
  wire wr_2841;
  wire wr_2842;
  wire wr_2843;
  wire wr_2844;
  wire wr_2845;
  wire wr_2846;
  wire wr_2847;
  wire wr_2848;
  wire wr_2849;
  wire wr_2850;
  wire wr_2851;
  wire wr_2852;
  wire wr_2853;
  wire wr_2854;
  wire wr_2855;
  wire wr_2856;
  wire wr_2857;
  wire wr_2858;
  wire wr_2859;
  wire wr_2860;
  wire wr_2861;
  wire wr_2862;
  wire wr_2863;
  wire wr_2864;
  wire wr_2865;
  wire wr_2866;
  wire wr_2867;
  wire wr_2868;
  wire wr_2869;
  wire wr_2870;
  wire wr_2871;
  wire wr_2872;
  wire wr_2873;
  wire wr_2874;
  wire wr_2875;
  wire wr_2876;
  wire wr_2877;
  wire wr_2878;
  wire wr_2879;
  wire wr_2880;
  wire wr_2881;
  wire wr_2882;
  wire wr_2883;
  wire wr_2884;
  wire wr_2885;
  wire wr_2886;
  wire wr_2887;
  wire wr_2888;
  wire wr_2889;
  wire wr_2890;
  wire wr_2891;
  wire wr_2892;
  wire wr_2893;
  wire wr_2894;
  wire wr_2895;
  wire wr_2896;
  wire wr_2897;
  wire wr_2898;
  wire wr_2899;
  wire wr_2900;
  wire wr_2901;
  wire wr_2902;
  wire wr_2903;
  wire wr_2904;
  wire wr_2905;
  wire wr_2906;
  wire wr_2907;
  wire wr_2908;
  wire wr_2909;
  wire wr_2910;

  not    g1( G599    ,           G348    );
  not    g2( G600    ,           G366    );
  not    g3( G612    ,           G358    );
  not    g4( wr_202  ,           G523    );
  not    g5( wr_203  ,           G341    );
  not    g6( wr_218  ,           G534    );
  not    g7( wr_219  ,           G351    );
  not    g8( wr_235  ,           G324    );
  not    g9( wr_250  ,           G514    );
  not   g10( wr_262  ,           G361    );
  not   g11( wr_267  ,           G479    );
  not   g12( wr_268  ,           G308    );
  not   g13( wr_285  ,           G490    );
  not   g14( wr_286  ,           G316    );
  not   g15( wr_306  ,           G302    );
  not   g16( wr_318  ,           G411    );
  not   g17( wr_319  ,           G273    );
  not   g18( wr_334  ,           G374    );
  not   g19( wr_335  ,           G281    );
  not   g20( wr_350  ,           G389    );
  not   g21( wr_351  ,           G257    );
  not   g22( wr_366  ,           G400    );
  not   g23( wr_367  ,           G265    );
  not   g24( wr_404  ,           G422    );
  not   g25( wr_405  ,           G226    );
  not   g26( wr_436  ,           G457    );
  not   g27( wr_437  ,           G210    );
  not   g28( wr_452  ,           G468    );
  not   g29( wr_453  ,           G218    );
  not   g30( wr_477  ,           G225    );
  not   g31( wr_478  ,           G335    );
  not   g32( wr_486  ,           G233    );
  not   g33( wr_502  ,           G217    );
  not   g34( wr_516  ,           G280    );
  not   g35( wr_524  ,           G288    );
  not   g36( wr_532  ,           G272    );
  not   g37( wr_548  ,           G264    );
  not   g38( wr_564  ,           G323    );
  not   g39( wr_565  ,           G332    );
  not   g40( wr_573  ,           G307    );
  not   g41( wr_582  ,           G315    );
  not   g42( wr_619  ,           G331    );
  not   g43( wr_421  ,           G234    );
  not   g44( wr_540  ,           G241    );
  not   g45( wr_234  ,           G503    );
  not   g46( wr_420  ,           G435    );
  not   g47( wr_389  ,           G206    );
  not   g48( wr_494  ,           G209    );
  not   g49( G593    ,           G299    );
  not   g50( wr_301  ,           G293    );
  not   g51( wr_261  ,           G248    );
  not   g52( wr_279  ,           G242    );
  not   g53( wr_388  ,           G446    );
  not   g54( wr_264  ,           G251    );
  not   g55( wr_277  ,           G254    );
  nor   g56( wr_2425 , G514    , G242    );
  not   g57( wr_863  ,           G54     );
  not   g58( wr_2252 ,           G2174   );
  not   g59( wr_723  ,           G289    );
  not   g60( wr_900  ,           G4      );
  not   g61( wr_1259 ,           G292    );
  not   g62( wr_677  ,           G369    );
  not   g63( wr_2526 ,           G1497   );
  not   g64( wr_1205 ,           G372    );
  nor   g65( wr_212  , G3548   , G341    );
  nor   g66( wr_228  , G3548   , G351    );
  nor   g67( wr_244  , G3548   , G324    );
  not   g68( wr_252  ,           G3546   );
  nor   g69( wr_328  , G3548   , G273    );
  nor   g70( wr_344  , G3548   , G281    );
  nor   g71( wr_360  , G3548   , G257    );
  nor   g72( wr_376  , G3548   , G265    );
  nor   g73( wr_414  , G3548   , G226    );
  nor   g74( wr_430  , G3548   , G234    );
  nor   g75( wr_446  , G3548   , G210    );
  nor   g76( wr_462  , G3548   , G218    );
  not   g77( wr_869  ,           G131    );
  not   g78( wr_870  ,           G4092   );
  not   g79( wr_889  ,           G129    );
  not   g80( wr_995  ,           G52     );
  not   g81( wr_1027 ,           G130    );
  not   g82( wr_1051 ,           G119    );
  not   g83( wr_1788 ,           G123    );
  not   g84( wr_1815 ,           G121    );
  not   g85( wr_1828 ,           G116    );
  not   g86( wr_1841 ,           G112    );
  not   g87( wr_861  ,           G4091   );
  not   g88( wr_907  ,           G117    );
  not   g89( wr_1108 ,           G122    );
  not   g90( wr_1140 ,           G128    );
  not   g91( wr_1164 ,           G127    );
  not   g92( wr_1184 ,           G126    );
  not   g93( wr_1870 ,           G115    );
  not   g94( wr_1883 ,           G114    );
  not   g95( wr_1896 ,           G53     );
  not   g96( wr_1909 ,           G113    );
  not   g97( wr_1450 ,           G1690   );
  not   g98( wr_1470 ,           G1694   );
  not   g99( wr_2837 ,           G94     );
  not  g100( wr_2879 ,           G179    );
  not  g101( wr_2883 ,           G176    );
  not  g102( G849    ,           G552    );
  not  g103( wr_129  ,           G27     );
  not  g104( wr_132  ,           G556    );
  not  g105( wr_135  ,           G31     );
  not  g106( wr_953  ,           G61     );
  not  g107( wr_954  ,           G4087   );
  not  g108( wr_958  ,           G11     );
  not  g109( wr_1068 ,           G4090   );
  not  g110( wr_1449 ,           G185    );
  not  g111( wr_1454 ,           G182    );
  not  g112( wr_1488 ,           G37     );
  not  g113( wr_1492 ,           G43     );
  not  g114( wr_1507 ,           G20     );
  not  g115( wr_1511 ,           G76     );
  not  g116( wr_1526 ,           G17     );
  not  g117( wr_1530 ,           G73     );
  not  g118( wr_1545 ,           G70     );
  not  g119( wr_1549 ,           G67     );
  not  g120( wr_1632 ,           G170    );
  not  g121( wr_1636 ,           G200    );
  not  g122( wr_1651 ,           G158    );
  not  g123( wr_1655 ,           G188    );
  not  g124( wr_1670 ,           G152    );
  not  g125( wr_1674 ,           G155    );
  not  g126( wr_1689 ,           G146    );
  not  g127( wr_1693 ,           G149    );
  not  g128( wr_1784 ,           G3717   );
  not  g129( wr_1925 ,           G106    );
  not  g130( wr_1929 ,           G109    );
  not  g131( wr_1961 ,           G49     );
  not  g132( wr_1965 ,           G46     );
  not  g133( wr_1980 ,           G103    );
  not  g134( wr_1984 ,           G100    );
  not  g135( wr_1999 ,           G40     );
  not  g136( wr_2003 ,           G91     );
  not  g137( wr_2069 ,           G173    );
  not  g138( wr_2073 ,           G203    );
  not  g139( wr_2088 ,           G167    );
  not  g140( wr_2092 ,           G197    );
  not  g141( wr_2107 ,           G164    );
  not  g142( wr_2111 ,           G194    );
  not  g143( wr_2126 ,           G161    );
  not  g144( wr_2130 ,           G191    );
  not  g145( wr_2472 ,           G120    );
  not  g146( wr_2812 ,           G118    );
  not  g147( wr_2843 ,           G64     );
  not  g148( wr_2847 ,           G14     );
  not  g149( wr_1442 ,           G1689   );
  not  g150( wr_1463 ,           G1691   );
  not  g151( wr_2826 ,           G97     );
  not  g152( wr_131  ,           G386    );
  not  g153( wr_160  ,           G24     );
  not  g154( wr_173  ,           G26     );
  not  g155( wr_184  ,           G79     );
  not  g156( wr_195  ,           G82     );
  not  g157( wr_946  ,           G4088   );
  not  g158( wr_1061 ,           G4089   );
  not  g159( wr_1773 ,           G3724   );
  not  g160( wr_1775 ,           G132    );
  not  g161( G850    ,           G562    );
  not  g162( G851    ,           G559    );
  not  g163( wr_156  ,           G25     );
  not  g164( wr_169  ,           G81     );
  not  g165( wr_180  ,           G23     );
  not  g166( wr_191  ,           G80     );
  not  g167( wr_138  ,           G87     );
  not  g168( wr_139  ,           G2358   );
  not  g169( wr_141  ,           G86     );
  not  g170( wr_145  ,           G34     );
  not  g171( wr_147  ,           G88     );
  not  g172( wr_151  ,           G83     );
  not  g173( G848    ,           G245    );
  not  g174( wr_134  ,           G140    );
  not  g175( wr_1441 ,           G137    );
  not  g176( wr_1770 ,           G135    );
  not  g177( wr_1771 ,           G4115   );
  not  g178( wr_124  ,           G141    );
  not  g179( wr_125  ,           G145    );
  not  g180( wr_126  ,           G1      );
  not  g181( wr_127  ,           G373    );
  not  g182( wr_128  ,           G136    );
  not  g183( G594    ,           G545    );
  not  g184( G602    ,           G549    );
  not  g185( G611    ,           G338    );
  not  g186( G144    ,           G141    );
  not  g187( G298    ,           G293    );
  not  g188( G973    ,           G3173   );
  not  g189( G603    ,           G545    );
  not  g190( G604    ,           G545    );
  not  g191( G926    ,           G137    );
  not  g192( G923    ,           G141    );
  not  g193( G921    ,           G1      );
  not  g194( G892    ,           G549    );
  not  g195( G887    ,           G299    );
  not  g196( G606    ,           G549    );
  not  g197( G993    ,           G1      );
  not  g198( G978    ,           G1      );
  not  g199( G949    ,           G1      );
  not  g200( G939    ,           G1      );
  not  g201( G889    ,           G299    );
  nor  g202( wr_476  , G335    , wr_453  );
  nor  g203( wr_479  , wr_478  , wr_477  );
  nor  g204( wr_485  , G335    , wr_405  );
  nor  g205( wr_487  , wr_478  , wr_486  );
  nor  g206( wr_501  , G335    , wr_437  );
  nor  g207( wr_503  , wr_478  , wr_502  );
  nor  g208( wr_515  , G335    , wr_319  );
  nor  g209( wr_517  , wr_478  , wr_516  );
  nor  g210( wr_523  , G335    , wr_335  );
  nor  g211( wr_525  , wr_478  , wr_524  );
  nor  g212( wr_531  , G335    , wr_367  );
  nor  g213( wr_533  , wr_478  , wr_532  );
  nor  g214( wr_547  , G335    , wr_351  );
  nor  g215( wr_549  , wr_478  , wr_548  );
  nor  g216( wr_563  , G332    , wr_286  );
  nor  g217( wr_566  , wr_565  , wr_564  );
  nor  g218( wr_572  , G332    , wr_306  );
  nor  g219( wr_574  , wr_565  , wr_573  );
  nor  g220( wr_581  , G332    , wr_268  );
  nor  g221( wr_583  , wr_565  , wr_582  );
  nor  g222( wr_595  , wr_262  , G332    );
  nor  g223( wr_596  , G600    , wr_565  );
  nor  g224( wr_599  , G338    , wr_565  );
  nor  g225( wr_604  , wr_203  , G332    );
  nor  g226( wr_605  , G599    , wr_565  );
  nor  g227( wr_611  , wr_219  , G332    );
  nor  g228( wr_612  , G612    , wr_565  );
  nor  g229( wr_618  , G332    , wr_235  );
  nor  g230( wr_620  , wr_565  , wr_619  );
  nor  g231( wr_539  , G335    , wr_421  );
  nor  g232( wr_541  , wr_478  , wr_540  );
  nor  g233( wr_493  , G335    , wr_389  );
  nor  g234( wr_495  , wr_478  , wr_494  );
  nor  g235( wr_577  , G332    , wr_301  );
  nor  g236( wr_578  , wr_565  , G593    );
  nor  g237( wr_207  , wr_202  , G341    );
  nor  g238( wr_223  , wr_218  , G351    );
  nor  g239( wr_239  , wr_234  , G324    );
  nor  g240( wr_2394 , wr_219  , wr_261  );
  nor  g241( wr_2407 , wr_203  , wr_261  );
  nor  g242( wr_2428 , wr_235  , wr_261  );
  nor  g243( wr_2401 , wr_219  , wr_279  );
  nor  g244( wr_2414 , wr_203  , wr_279  );
  nor  g245( wr_2435 , wr_235  , wr_279  );
  nor  g246( wr_323  , wr_318  , G273    );
  nor  g247( wr_355  , wr_350  , G257    );
  nor  g248( wr_371  , wr_366  , G265    );
  nor  g249( wr_425  , wr_420  , G234    );
  nor  g250( wr_2713 , wr_319  , wr_261  );
  nor  g251( wr_2726 , wr_367  , wr_261  );
  nor  g252( wr_2743 , wr_351  , wr_261  );
  nor  g253( wr_2756 , wr_261  , wr_421  );
  nor  g254( wr_2400 , G351    , wr_277  );
  nor  g255( wr_2413 , G341    , wr_277  );
  nor  g256( wr_2434 , G324    , wr_277  );
  nor  g257( wr_2720 , wr_319  , wr_279  );
  nor  g258( wr_2733 , wr_367  , wr_279  );
  nor  g259( wr_2750 , wr_351  , wr_279  );
  nor  g260( wr_2763 , wr_279  , wr_421  );
  nor  g261( wr_269  , wr_268  , wr_261  );
  nor  g262( wr_272  , wr_267  , G308    );
  nor  g263( wr_287  , wr_286  , wr_261  );
  nor  g264( wr_290  , wr_285  , G316    );
  nor  g265( wr_2424 , wr_250  , wr_261  );
  nor  g266( wr_280  , wr_268  , wr_279  );
  nor  g267( wr_296  , wr_286  , wr_279  );
  nor  g268( wr_339  , wr_334  , G281    );
  nor  g269( wr_2719 , G273    , wr_277  );
  nor  g270( wr_2732 , G265    , wr_277  );
  nor  g271( wr_2749 , G257    , wr_277  );
  nor  g272( wr_2762 , wr_277  , G234    );
  nor  g273( wr_2773 , wr_335  , wr_261  );
  nor  g274( wr_390  , wr_261  , wr_389  );
  nor  g275( wr_393  , wr_388  , G206    );
  nor  g276( wr_409  , wr_404  , G226    );
  nor  g277( wr_441  , wr_436  , G210    );
  nor  g278( wr_457  , wr_452  , G218    );
  nor  g279( wr_2663 , wr_261  , wr_405  );
  nor  g280( wr_2676 , wr_261  , wr_453  );
  nor  g281( wr_2692 , wr_261  , wr_437  );
  nor  g282( wr_2780 , wr_335  , wr_279  );
  nor  g283( wr_263  , wr_262  , wr_261  );
  nor  g284( wr_265  , G361    , wr_264  );
  nor  g285( wr_278  , G308    , wr_277  );
  nor  g286( wr_295  , G316    , wr_277  );
  nor  g287( wr_399  , wr_279  , wr_389  );
  nor  g288( wr_2670 , wr_279  , wr_405  );
  nor  g289( wr_2683 , wr_279  , wr_453  );
  nor  g290( wr_2699 , wr_279  , wr_437  );
  nor  g291( wr_302  , wr_301  , wr_279  );
  nor  g292( wr_303  , G293    , wr_277  );
  nor  g293( wr_307  , wr_306  , wr_261  );
  nor  g294( wr_308  , G302    , wr_264  );
  nor  g295( wr_1258 , G335    , wr_723  );
  nor  g296( wr_1260 , wr_478  , wr_1259 );
  nor  g297( wr_2779 , G281    , wr_277  );
  nor  g298( wr_398  , wr_277  , G206    );
  nor  g299( wr_673  , wr_219  , G341    );
  nor  g300( wr_674  , G351    , wr_203  );
  nor  g301( wr_678  , wr_677  , G361    );
  nor  g302( wr_679  , G369    , wr_262  );
  nor  g303( wr_715  , wr_319  , G265    );
  nor  g304( wr_716  , G273    , wr_367  );
  nor  g305( wr_719  , wr_351  , G234    );
  nor  g306( wr_720  , G257    , wr_421  );
  nor  g307( wr_724  , wr_723  , G281    );
  nor  g308( wr_725  , G289    , wr_335  );
  nor  g309( wr_2669 , wr_277  , G226    );
  nor  g310( wr_2682 , wr_277  , G218    );
  nor  g311( wr_2698 , wr_277  , G210    );
  nor  g312( wr_204  , G3552   , wr_203  );
  nor  g313( wr_220  , G3552   , wr_219  );
  nor  g314( wr_236  , G3552   , wr_235  );
  nor  g315( wr_213  , G3546   , wr_203  );
  nor  g316( wr_229  , G3546   , wr_219  );
  nor  g317( wr_245  , G3546   , wr_235  );
  nor  g318( wr_1204 , wr_677  , G332    );
  nor  g319( wr_1206 , wr_1205 , wr_565  );
  nor  g320( wr_320  , G3552   , wr_319  );
  nor  g321( wr_336  , G3552   , wr_335  );
  nor  g322( wr_352  , G3552   , wr_351  );
  nor  g323( wr_368  , G3552   , wr_367  );
  nor  g324( wr_406  , G3552   , wr_405  );
  nor  g325( wr_422  , G3552   , wr_421  );
  nor  g326( wr_438  , G3552   , wr_437  );
  nor  g327( wr_454  , G3552   , wr_453  );
  nor  g328( wr_662  , wr_286  , G308    );
  nor  g329( wr_663  , G316    , wr_268  );
  nor  g330( wr_665  , wr_306  , G293    );
  nor  g331( wr_666  , G302    , wr_301  );
  nor  g332( wr_704  , wr_405  , G218    );
  nor  g333( wr_705  , G226    , wr_453  );
  nor  g334( wr_707  , wr_437  , G206    );
  nor  g335( wr_708  , G210    , wr_389  );
  nor  g336( wr_329  , G3546   , wr_319  );
  nor  g337( wr_345  , G3546   , wr_335  );
  nor  g338( wr_361  , G3546   , wr_351  );
  nor  g339( wr_377  , G3546   , wr_367  );
  nor  g340( wr_415  , G3546   , wr_405  );
  nor  g341( wr_431  , G3546   , wr_421  );
  nor  g342( wr_447  , G3546   , wr_437  );
  nor  g343( wr_463  , G3546   , wr_453  );
  nor  g344( wr_251  , G3552   , wr_250  );
  nor  g345( wr_253  , wr_252  , G514    );
  nor  g346( wr_871  , wr_870  , wr_869  );
  nor  g347( wr_890  , wr_870  , wr_889  );
  nor  g348( wr_996  , wr_870  , wr_995  );
  nor  g349( wr_1028 , wr_870  , wr_1027 );
  nor  g350( wr_1052 , wr_870  , wr_1051 );
  nor  g351( wr_1804 , wr_870  , wr_1788 );
  nor  g352( wr_1816 , wr_870  , wr_1815 );
  nor  g353( wr_1829 , wr_870  , wr_1828 );
  nor  g354( wr_1842 , wr_870  , wr_1841 );
  nor  g355( wr_908  , wr_870  , wr_907  );
  nor  g356( wr_1109 , wr_870  , wr_1108 );
  nor  g357( wr_1141 , wr_870  , wr_1140 );
  nor  g358( wr_1165 , wr_870  , wr_1164 );
  nor  g359( wr_1185 , wr_870  , wr_1184 );
  nor  g360( wr_1871 , wr_870  , wr_1870 );
  nor  g361( wr_1884 , wr_870  , wr_1883 );
  nor  g362( wr_1897 , wr_870  , wr_1896 );
  nor  g363( wr_1910 , wr_870  , wr_1909 );
  nor  g364( wr_2838 , wr_870  , wr_2837 );
  nor  g365( wr_2880 , wr_1450 , wr_2879 );
  nor  g366( wr_2884 , wr_1450 , wr_2883 );
  nor  g367( wr_2899 , wr_1470 , wr_2879 );
  nor  g368( wr_2902 , wr_1470 , wr_2883 );
  nor  g369( wr_136  , wr_135  , wr_129  );
  nor  g370( wr_955  , wr_954  , wr_953  );
  nor  g371( wr_959  , wr_954  , wr_958  );
  nor  g372( wr_1069 , wr_1068 , wr_953  );
  nor  g373( wr_1072 , wr_1068 , wr_958  );
  nor  g374( wr_1451 , wr_1450 , wr_1449 );
  nor  g375( wr_1455 , wr_1450 , wr_1454 );
  nor  g376( wr_1471 , wr_1470 , wr_1449 );
  nor  g377( wr_1474 , wr_1470 , wr_1454 );
  nor  g378( wr_1489 , wr_954  , wr_1488 );
  nor  g379( wr_1493 , wr_954  , wr_1492 );
  nor  g380( wr_1508 , wr_954  , wr_1507 );
  nor  g381( wr_1512 , wr_954  , wr_1511 );
  nor  g382( wr_1527 , wr_954  , wr_1526 );
  nor  g383( wr_1531 , wr_954  , wr_1530 );
  nor  g384( wr_1546 , wr_954  , wr_1545 );
  nor  g385( wr_1550 , wr_954  , wr_1549 );
  nor  g386( wr_1564 , wr_1068 , wr_1488 );
  nor  g387( wr_1567 , wr_1068 , wr_1492 );
  nor  g388( wr_1581 , wr_1068 , wr_1507 );
  nor  g389( wr_1584 , wr_1068 , wr_1511 );
  nor  g390( wr_1598 , wr_1068 , wr_1526 );
  nor  g391( wr_1601 , wr_1068 , wr_1530 );
  nor  g392( wr_1615 , wr_1068 , wr_1545 );
  nor  g393( wr_1618 , wr_1068 , wr_1549 );
  nor  g394( wr_1633 , wr_1450 , wr_1632 );
  nor  g395( wr_1637 , wr_1450 , wr_1636 );
  nor  g396( wr_1652 , wr_1450 , wr_1651 );
  nor  g397( wr_1656 , wr_1450 , wr_1655 );
  nor  g398( wr_1671 , wr_1450 , wr_1670 );
  nor  g399( wr_1675 , wr_1450 , wr_1674 );
  nor  g400( wr_1690 , wr_1450 , wr_1689 );
  nor  g401( wr_1694 , wr_1450 , wr_1693 );
  nor  g402( wr_1708 , wr_1470 , wr_1632 );
  nor  g403( wr_1711 , wr_1470 , wr_1636 );
  nor  g404( wr_1725 , wr_1470 , wr_1651 );
  nor  g405( wr_1728 , wr_1470 , wr_1655 );
  nor  g406( wr_1742 , wr_1470 , wr_1670 );
  nor  g407( wr_1745 , wr_1470 , wr_1674 );
  nor  g408( wr_1759 , wr_1470 , wr_1689 );
  nor  g409( wr_1762 , wr_1470 , wr_1693 );
  nor  g410( wr_1789 , wr_1784 , wr_1788 );
  nor  g411( wr_1859 , wr_132  , G849    );
  nor  g412( wr_1926 , wr_1068 , wr_1925 );
  nor  g413( wr_1930 , wr_1068 , wr_1929 );
  nor  g414( wr_1944 , wr_954  , wr_1925 );
  nor  g415( wr_1947 , wr_954  , wr_1929 );
  nor  g416( wr_1962 , wr_954  , wr_1961 );
  nor  g417( wr_1966 , wr_954  , wr_1965 );
  nor  g418( wr_1981 , wr_954  , wr_1980 );
  nor  g419( wr_1985 , wr_954  , wr_1984 );
  nor  g420( wr_2000 , wr_954  , wr_1999 );
  nor  g421( wr_2004 , wr_954  , wr_2003 );
  nor  g422( wr_2018 , wr_1068 , wr_1961 );
  nor  g423( wr_2021 , wr_1068 , wr_1965 );
  nor  g424( wr_2035 , wr_1068 , wr_1980 );
  nor  g425( wr_2038 , wr_1068 , wr_1984 );
  nor  g426( wr_2052 , wr_1068 , wr_1999 );
  nor  g427( wr_2055 , wr_1068 , wr_2003 );
  nor  g428( wr_2070 , wr_1450 , wr_2069 );
  nor  g429( wr_2074 , wr_1450 , wr_2073 );
  nor  g430( wr_2089 , wr_1450 , wr_2088 );
  nor  g431( wr_2093 , wr_1450 , wr_2092 );
  nor  g432( wr_2108 , wr_1450 , wr_2107 );
  nor  g433( wr_2112 , wr_1450 , wr_2111 );
  nor  g434( wr_2127 , wr_1450 , wr_2126 );
  nor  g435( wr_2131 , wr_1450 , wr_2130 );
  nor  g436( wr_2145 , wr_1470 , wr_2069 );
  nor  g437( wr_2148 , wr_1470 , wr_2073 );
  nor  g438( wr_2162 , wr_1470 , wr_2088 );
  nor  g439( wr_2165 , wr_1470 , wr_2092 );
  nor  g440( wr_2179 , wr_1470 , wr_2107 );
  nor  g441( wr_2182 , wr_1470 , wr_2111 );
  nor  g442( wr_2196 , wr_1470 , wr_2126 );
  nor  g443( wr_2199 , wr_1470 , wr_2130 );
  nor  g444( wr_2473 , wr_870  , wr_2472 );
  nor  g445( wr_2813 , wr_870  , wr_2812 );
  nor  g446( wr_2844 , wr_954  , wr_2843 );
  nor  g447( wr_2848 , wr_954  , wr_2847 );
  nor  g448( wr_2862 , wr_1068 , wr_2843 );
  nor  g449( wr_2865 , wr_1068 , wr_2847 );
  nor  g450( wr_2827 , wr_870  , wr_2826 );
  nor  g451( wr_2471 , wr_870  , wr_861  );
  nor  g452( wr_164  , wr_135  , wr_129  );
  nor  g453( wr_140  , wr_139  , wr_138  );
  nor  g454( wr_142  , G2358   , wr_141  );
  nor  g455( wr_146  , wr_139  , wr_145  );
  nor  g456( wr_148  , G2358   , wr_147  );
  nor  g457( wr_152  , wr_139  , wr_151  );
  nor  g458( wr_153  , G2358   , wr_151  );
  nor  g459( wr_130  , G2824   , wr_129  );
  nor  g460( wr_133  , wr_132  , wr_131  );
  nor  g461( wr_1772 , wr_1771 , wr_1770 );
  nor  g462( G601    , G850    , G849    );
  nor  g463( G810    , wr_125  , wr_124  );
  nor  g464( G634    , wr_127  , wr_126  );
  nor  g465( G815    , G3173   , wr_128  );
  nor  g466( wr_480  , wr_479  , wr_476  );
  nor  g467( wr_488  , wr_487  , wr_485  );
  nor  g468( wr_504  , wr_503  , wr_501  );
  nor  g469( wr_518  , wr_517  , wr_515  );
  nor  g470( wr_526  , wr_525  , wr_523  );
  nor  g471( wr_534  , wr_533  , wr_531  );
  nor  g472( wr_550  , wr_549  , wr_547  );
  nor  g473( wr_567  , wr_566  , wr_563  );
  nor  g474( wr_575  , wr_574  , wr_572  );
  nor  g475( wr_584  , wr_583  , wr_581  );
  nor  g476( wr_597  , wr_596  , wr_595  );
  not  g477( wr_600  ,           wr_599  );
  nor  g478( wr_602  , wr_599  , G514    );
  nor  g479( wr_606  , wr_605  , wr_604  );
  nor  g480( wr_613  , wr_612  , wr_611  );
  nor  g481( wr_621  , wr_620  , wr_618  );
  nor  g482( wr_825  , wr_599  , wr_250  );
  nor  g483( wr_542  , wr_541  , wr_539  );
  nor  g484( wr_496  , wr_495  , wr_493  );
  nor  g485( wr_579  , wr_578  , wr_577  );
  not  g486( wr_208  ,           wr_207  );
  not  g487( wr_224  ,           wr_223  );
  not  g488( wr_240  ,           wr_239  );
  not  g489( wr_2395 ,           wr_2394 );
  not  g490( wr_2408 ,           wr_2407 );
  not  g491( wr_2429 ,           wr_2428 );
  nor  g492( wr_2402 , wr_2401 , G534    );
  nor  g493( wr_2415 , wr_2414 , G523    );
  nor  g494( wr_2436 , wr_2435 , G503    );
  not  g495( wr_324  ,           wr_323  );
  not  g496( wr_356  ,           wr_355  );
  not  g497( wr_372  ,           wr_371  );
  not  g498( wr_426  ,           wr_425  );
  not  g499( wr_2714 ,           wr_2713 );
  not  g500( wr_2727 ,           wr_2726 );
  not  g501( wr_2744 ,           wr_2743 );
  not  g502( wr_2757 ,           wr_2756 );
  nor  g503( wr_2721 , wr_2720 , G411    );
  nor  g504( wr_2734 , wr_2733 , G400    );
  nor  g505( wr_2751 , wr_2750 , G389    );
  nor  g506( wr_2764 , wr_2763 , G435    );
  not  g507( wr_270  ,           wr_269  );
  not  g508( wr_273  ,           wr_272  );
  not  g509( wr_288  ,           wr_287  );
  not  g510( wr_291  ,           wr_290  );
  nor  g511( wr_2426 , wr_2425 , wr_2424 );
  nor  g512( wr_281  , wr_280  , G479    );
  nor  g513( wr_297  , wr_296  , G490    );
  not  g514( wr_340  ,           wr_339  );
  not  g515( wr_2774 ,           wr_2773 );
  not  g516( wr_391  ,           wr_390  );
  not  g517( wr_394  ,           wr_393  );
  not  g518( wr_410  ,           wr_409  );
  not  g519( wr_442  ,           wr_441  );
  not  g520( wr_458  ,           wr_457  );
  not  g521( wr_2664 ,           wr_2663 );
  not  g522( wr_2677 ,           wr_2676 );
  not  g523( wr_2693 ,           wr_2692 );
  nor  g524( wr_2781 , wr_2780 , G374    );
  nor  g525( wr_266  , wr_265  , wr_263  );
  nor  g526( wr_400  , wr_399  , G446    );
  nor  g527( wr_2671 , wr_2670 , G422    );
  nor  g528( wr_2684 , wr_2683 , G468    );
  nor  g529( wr_2700 , wr_2699 , G457    );
  nor  g530( wr_304  , wr_303  , wr_302  );
  nor  g531( wr_309  , wr_308  , wr_307  );
  nor  g532( wr_1261 , wr_1260 , wr_1258 );
  nor  g533( wr_675  , wr_674  , wr_673  );
  nor  g534( wr_680  , wr_679  , wr_678  );
  nor  g535( wr_717  , wr_716  , wr_715  );
  nor  g536( wr_721  , wr_720  , wr_719  );
  nor  g537( wr_726  , wr_725  , wr_724  );
  not  g538( wr_205  ,           wr_204  );
  not  g539( wr_221  ,           wr_220  );
  not  g540( wr_237  ,           wr_236  );
  nor  g541( wr_214  , wr_213  , G523    );
  nor  g542( wr_230  , wr_229  , G534    );
  nor  g543( wr_246  , wr_245  , G503    );
  nor  g544( wr_1207 , wr_1206 , wr_1204 );
  not  g545( wr_321  ,           wr_320  );
  not  g546( wr_337  ,           wr_336  );
  not  g547( wr_353  ,           wr_352  );
  not  g548( wr_369  ,           wr_368  );
  not  g549( wr_407  ,           wr_406  );
  not  g550( wr_423  ,           wr_422  );
  not  g551( wr_439  ,           wr_438  );
  not  g552( wr_455  ,           wr_454  );
  nor  g553( wr_664  , wr_663  , wr_662  );
  nor  g554( wr_667  , wr_666  , wr_665  );
  nor  g555( wr_706  , wr_705  , wr_704  );
  nor  g556( wr_709  , wr_708  , wr_707  );
  nor  g557( wr_330  , wr_329  , G411    );
  nor  g558( wr_346  , wr_345  , G374    );
  nor  g559( wr_362  , wr_361  , G389    );
  nor  g560( wr_378  , wr_377  , G400    );
  nor  g561( wr_416  , wr_415  , G422    );
  nor  g562( wr_432  , wr_431  , G435    );
  nor  g563( wr_448  , wr_447  , G457    );
  nor  g564( wr_464  , wr_463  , G468    );
  nor  g565( wr_254  , wr_253  , wr_251  );
  not  g566( wr_872  ,           wr_871  );
  not  g567( wr_891  ,           wr_890  );
  not  g568( wr_997  ,           wr_996  );
  not  g569( wr_1029 ,           wr_1028 );
  not  g570( wr_1053 ,           wr_1052 );
  not  g571( wr_1805 ,           wr_1804 );
  not  g572( wr_1817 ,           wr_1816 );
  not  g573( wr_1830 ,           wr_1829 );
  not  g574( wr_1843 ,           wr_1842 );
  not  g575( wr_909  ,           wr_908  );
  not  g576( wr_1110 ,           wr_1109 );
  not  g577( wr_1142 ,           wr_1141 );
  not  g578( wr_1166 ,           wr_1165 );
  not  g579( wr_1186 ,           wr_1185 );
  not  g580( wr_1872 ,           wr_1871 );
  not  g581( wr_1885 ,           wr_1884 );
  not  g582( wr_1898 ,           wr_1897 );
  not  g583( wr_1911 ,           wr_1910 );
  not  g584( wr_2881 ,           wr_2880 );
  not  g585( wr_2885 ,           wr_2884 );
  not  g586( wr_2900 ,           wr_2899 );
  not  g587( wr_2903 ,           wr_2902 );
  not  g588( G809    ,           wr_136  );
  not  g589( wr_956  ,           wr_955  );
  not  g590( wr_960  ,           wr_959  );
  not  g591( wr_1070 ,           wr_1069 );
  not  g592( wr_1073 ,           wr_1072 );
  not  g593( wr_1452 ,           wr_1451 );
  not  g594( wr_1456 ,           wr_1455 );
  not  g595( wr_1472 ,           wr_1471 );
  not  g596( wr_1475 ,           wr_1474 );
  not  g597( wr_1490 ,           wr_1489 );
  not  g598( wr_1494 ,           wr_1493 );
  not  g599( wr_1509 ,           wr_1508 );
  not  g600( wr_1513 ,           wr_1512 );
  not  g601( wr_1528 ,           wr_1527 );
  not  g602( wr_1532 ,           wr_1531 );
  not  g603( wr_1547 ,           wr_1546 );
  not  g604( wr_1551 ,           wr_1550 );
  not  g605( wr_1565 ,           wr_1564 );
  not  g606( wr_1568 ,           wr_1567 );
  not  g607( wr_1582 ,           wr_1581 );
  not  g608( wr_1585 ,           wr_1584 );
  not  g609( wr_1599 ,           wr_1598 );
  not  g610( wr_1602 ,           wr_1601 );
  not  g611( wr_1616 ,           wr_1615 );
  not  g612( wr_1619 ,           wr_1618 );
  not  g613( wr_1634 ,           wr_1633 );
  not  g614( wr_1638 ,           wr_1637 );
  not  g615( wr_1653 ,           wr_1652 );
  not  g616( wr_1657 ,           wr_1656 );
  not  g617( wr_1672 ,           wr_1671 );
  not  g618( wr_1676 ,           wr_1675 );
  not  g619( wr_1691 ,           wr_1690 );
  not  g620( wr_1695 ,           wr_1694 );
  not  g621( wr_1709 ,           wr_1708 );
  not  g622( wr_1712 ,           wr_1711 );
  not  g623( wr_1726 ,           wr_1725 );
  not  g624( wr_1729 ,           wr_1728 );
  not  g625( wr_1743 ,           wr_1742 );
  not  g626( wr_1746 ,           wr_1745 );
  not  g627( wr_1760 ,           wr_1759 );
  not  g628( wr_1763 ,           wr_1762 );
  not  g629( wr_1790 ,           wr_1789 );
  not  g630( wr_1860 ,           wr_1859 );
  not  g631( wr_1927 ,           wr_1926 );
  not  g632( wr_1931 ,           wr_1930 );
  not  g633( wr_1945 ,           wr_1944 );
  not  g634( wr_1948 ,           wr_1947 );
  not  g635( wr_1963 ,           wr_1962 );
  not  g636( wr_1967 ,           wr_1966 );
  not  g637( wr_1982 ,           wr_1981 );
  not  g638( wr_1986 ,           wr_1985 );
  not  g639( wr_2001 ,           wr_2000 );
  not  g640( wr_2005 ,           wr_2004 );
  not  g641( wr_2019 ,           wr_2018 );
  not  g642( wr_2022 ,           wr_2021 );
  not  g643( wr_2036 ,           wr_2035 );
  not  g644( wr_2039 ,           wr_2038 );
  not  g645( wr_2053 ,           wr_2052 );
  not  g646( wr_2056 ,           wr_2055 );
  not  g647( wr_2071 ,           wr_2070 );
  not  g648( wr_2075 ,           wr_2074 );
  not  g649( wr_2090 ,           wr_2089 );
  not  g650( wr_2094 ,           wr_2093 );
  not  g651( wr_2109 ,           wr_2108 );
  not  g652( wr_2113 ,           wr_2112 );
  not  g653( wr_2128 ,           wr_2127 );
  not  g654( wr_2132 ,           wr_2131 );
  not  g655( wr_2146 ,           wr_2145 );
  not  g656( wr_2149 ,           wr_2148 );
  not  g657( wr_2163 ,           wr_2162 );
  not  g658( wr_2166 ,           wr_2165 );
  not  g659( wr_2180 ,           wr_2179 );
  not  g660( wr_2183 ,           wr_2182 );
  not  g661( wr_2197 ,           wr_2196 );
  not  g662( wr_2200 ,           wr_2199 );
  not  g663( wr_2474 ,           wr_2473 );
  not  g664( wr_2814 ,           wr_2813 );
  not  g665( wr_2845 ,           wr_2844 );
  not  g666( wr_2849 ,           wr_2848 );
  not  g667( wr_2863 ,           wr_2862 );
  not  g668( wr_2866 ,           wr_2865 );
  not  g669( wr_165  ,           wr_164  );
  nor  g670( wr_143  , wr_142  , wr_140  );
  nor  g671( wr_149  , wr_148  , wr_146  );
  nor  g672( wr_154  , wr_153  , wr_152  );
  not  g673( G845    ,           wr_130  );
  not  g674( G847    ,           wr_133  );
  nor  g675( wr_481  , wr_480  , G468    );
  not  g676( wr_482  ,           wr_480  );
  nor  g677( wr_489  , wr_488  , G422    );
  not  g678( wr_490  ,           wr_488  );
  nor  g679( wr_505  , wr_504  , G457    );
  not  g680( wr_506  ,           wr_504  );
  nor  g681( wr_519  , wr_518  , G411    );
  not  g682( wr_520  ,           wr_518  );
  nor  g683( wr_527  , wr_526  , G374    );
  not  g684( wr_528  ,           wr_526  );
  nor  g685( wr_535  , wr_534  , G400    );
  not  g686( wr_536  ,           wr_534  );
  nor  g687( wr_551  , wr_550  , G389    );
  not  g688( wr_552  ,           wr_550  );
  not  g689( wr_568  ,           wr_567  );
  nor  g690( wr_570  , wr_567  , G490    );
  not  g691( wr_576  ,           wr_575  );
  not  g692( wr_585  ,           wr_584  );
  nor  g693( wr_587  , wr_584  , G479    );
  not  g694( wr_598  ,           wr_597  );
  nor  g695( wr_601  , wr_600  , wr_250  );
  not  g696( wr_607  ,           wr_606  );
  nor  g697( wr_609  , wr_606  , G523    );
  not  g698( wr_614  ,           wr_613  );
  nor  g699( wr_616  , wr_613  , G534    );
  nor  g700( wr_754  , wr_488  , wr_404  );
  nor  g701( wr_761  , wr_480  , wr_452  );
  nor  g702( wr_776  , wr_534  , wr_366  );
  nor  g703( wr_781  , wr_526  , wr_334  );
  nor  g704( wr_790  , wr_518  , wr_318  );
  nor  g705( wr_807  , wr_567  , wr_285  );
  nor  g706( wr_814  , wr_584  , wr_267  );
  nor  g707( wr_829  , wr_606  , wr_202  );
  nor  g708( wr_841  , wr_613  , wr_218  );
  nor  g709( wr_750  , wr_504  , wr_436  );
  not  g710( wr_622  ,           wr_621  );
  nor  g711( wr_624  , wr_621  , G503    );
  nor  g712( wr_772  , wr_550  , wr_350  );
  not  g713( wr_544  ,           wr_542  );
  nor  g714( wr_543  , wr_542  , G435    );
  not  g715( wr_498  ,           wr_496  );
  nor  g716( wr_497  , wr_496  , G446    );
  not  g717( wr_580  ,           wr_579  );
  nor  g718( wr_828  , wr_621  , wr_234  );
  nor  g719( wr_2396 , wr_2395 , wr_218  );
  nor  g720( wr_2397 , wr_224  , wr_264  );
  nor  g721( wr_2409 , wr_2408 , wr_202  );
  nor  g722( wr_2410 , wr_208  , wr_264  );
  nor  g723( wr_2430 , wr_2429 , wr_234  );
  nor  g724( wr_2431 , wr_240  , wr_264  );
  not  g725( wr_826  ,           wr_825  );
  not  g726( wr_2403 ,           wr_2402 );
  not  g727( wr_2416 ,           wr_2415 );
  not  g728( wr_2437 ,           wr_2436 );
  nor  g729( wr_775  , wr_542  , wr_420  );
  nor  g730( wr_2715 , wr_2714 , wr_318  );
  nor  g731( wr_2716 , wr_324  , wr_264  );
  nor  g732( wr_2728 , wr_2727 , wr_366  );
  nor  g733( wr_2729 , wr_372  , wr_264  );
  nor  g734( wr_2745 , wr_2744 , wr_350  );
  nor  g735( wr_2746 , wr_356  , wr_264  );
  nor  g736( wr_2758 , wr_2757 , wr_420  );
  nor  g737( wr_2759 , wr_426  , wr_264  );
  not  g738( wr_2722 ,           wr_2721 );
  not  g739( wr_2735 ,           wr_2734 );
  not  g740( wr_2752 ,           wr_2751 );
  not  g741( wr_2765 ,           wr_2764 );
  nor  g742( wr_271  , wr_270  , wr_267  );
  nor  g743( wr_274  , wr_273  , wr_264  );
  nor  g744( wr_289  , wr_288  , wr_285  );
  nor  g745( wr_292  , wr_291  , wr_264  );
  not  g746( wr_2427 ,           wr_2426 );
  not  g747( wr_282  ,           wr_281  );
  not  g748( wr_298  ,           wr_297  );
  nor  g749( wr_2775 , wr_2774 , wr_334  );
  nor  g750( wr_2776 , wr_340  , wr_264  );
  nor  g751( wr_392  , wr_391  , wr_388  );
  nor  g752( wr_395  , wr_394  , wr_264  );
  nor  g753( wr_2665 , wr_2664 , wr_404  );
  nor  g754( wr_2666 , wr_410  , wr_264  );
  nor  g755( wr_2678 , wr_2677 , wr_452  );
  nor  g756( wr_2679 , wr_458  , wr_264  );
  nor  g757( wr_2694 , wr_2693 , wr_436  );
  nor  g758( wr_2695 , wr_442  , wr_264  );
  not  g759( wr_2782 ,           wr_2781 );
  not  g760( wr_401  ,           wr_400  );
  not  g761( wr_874  ,           wr_266  );
  not  g762( wr_2672 ,           wr_2671 );
  not  g763( wr_2685 ,           wr_2684 );
  not  g764( wr_2701 ,           wr_2700 );
  not  g765( wr_305  ,           wr_304  );
  not  g766( wr_1262 ,           wr_1261 );
  not  g767( wr_1819 ,           wr_309  );
  not  g768( wr_676  ,           wr_675  );
  not  g769( wr_684  ,           wr_680  );
  not  g770( wr_718  ,           wr_717  );
  not  g771( wr_722  ,           wr_721  );
  not  g772( wr_730  ,           wr_726  );
  nor  g773( wr_2387 , wr_309  , wr_304  );
  nor  g774( wr_681  , wr_680  , wr_235  );
  nor  g775( wr_693  , wr_675  , G324    );
  nor  g776( wr_739  , wr_721  , wr_717  );
  nor  g777( wr_206  , wr_205  , wr_202  );
  nor  g778( wr_209  , wr_208  , G3550   );
  nor  g779( wr_222  , wr_221  , wr_218  );
  nor  g780( wr_225  , wr_224  , G3550   );
  nor  g781( wr_238  , wr_237  , wr_234  );
  nor  g782( wr_241  , wr_240  , G3550   );
  not  g783( wr_215  ,           wr_214  );
  not  g784( wr_231  ,           wr_230  );
  not  g785( wr_247  ,           wr_246  );
  not  g786( wr_1208 ,           wr_1207 );
  nor  g787( wr_322  , wr_321  , wr_318  );
  nor  g788( wr_325  , wr_324  , G3550   );
  nor  g789( wr_338  , wr_337  , wr_334  );
  nor  g790( wr_341  , wr_340  , G3550   );
  nor  g791( wr_354  , wr_353  , wr_350  );
  nor  g792( wr_357  , wr_356  , G3550   );
  nor  g793( wr_370  , wr_369  , wr_366  );
  nor  g794( wr_373  , wr_372  , G3550   );
  nor  g795( wr_408  , wr_407  , wr_404  );
  nor  g796( wr_411  , wr_410  , G3550   );
  nor  g797( wr_424  , wr_423  , wr_420  );
  nor  g798( wr_427  , wr_426  , G3550   );
  nor  g799( wr_440  , wr_439  , wr_436  );
  nor  g800( wr_443  , wr_442  , G3550   );
  nor  g801( wr_456  , wr_455  , wr_452  );
  nor  g802( wr_459  , wr_458  , G3550   );
  not  g803( wr_668  ,           wr_667  );
  not  g804( wr_670  ,           wr_664  );
  not  g805( wr_710  ,           wr_709  );
  not  g806( wr_712  ,           wr_706  );
  nor  g807( wr_1214 , wr_621  , wr_600  );
  not  g808( wr_331  ,           wr_330  );
  not  g809( wr_347  ,           wr_346  );
  not  g810( wr_363  ,           wr_362  );
  not  g811( wr_379  ,           wr_378  );
  not  g812( wr_417  ,           wr_416  );
  not  g813( wr_433  ,           wr_432  );
  not  g814( wr_449  ,           wr_448  );
  not  g815( wr_465  ,           wr_464  );
  not  g816( wr_1031 ,           wr_254  );
  nor  g817( wr_864  , wr_597  , wr_863  );
  nor  g818( wr_1807 , wr_304  , G4092   );
  nor  g819( wr_873  , wr_872  , G4091   );
  nor  g820( wr_892  , wr_891  , G4091   );
  nor  g821( wr_998  , wr_997  , G4091   );
  nor  g822( wr_1030 , wr_1029 , G4091   );
  nor  g823( wr_1054 , wr_1053 , G4091   );
  nor  g824( wr_1806 , wr_1805 , G4091   );
  nor  g825( wr_1818 , wr_1817 , G4091   );
  nor  g826( wr_1831 , wr_1830 , G4091   );
  nor  g827( wr_1844 , wr_1843 , G4091   );
  nor  g828( wr_910  , wr_909  , G4091   );
  nor  g829( wr_1111 , wr_1110 , G4091   );
  nor  g830( wr_1143 , wr_1142 , G4091   );
  nor  g831( wr_1167 , wr_1166 , G4091   );
  nor  g832( wr_1187 , wr_1186 , G4091   );
  nor  g833( wr_1873 , wr_1872 , G4091   );
  nor  g834( wr_1886 , wr_1885 , G4091   );
  nor  g835( wr_1899 , wr_1898 , G4091   );
  nor  g836( wr_1912 , wr_1911 , G4091   );
  nor  g837( wr_2882 , wr_2881 , wr_1442 );
  nor  g838( wr_2886 , wr_2885 , G1689   );
  nor  g839( wr_2901 , wr_2900 , wr_1463 );
  nor  g840( wr_2904 , wr_2903 , G1691   );
  nor  g841( wr_161  , G809    , wr_160  );
  nor  g842( wr_174  , G809    , wr_173  );
  nor  g843( wr_185  , G809    , wr_184  );
  nor  g844( wr_196  , G809    , wr_195  );
  nor  g845( wr_753  , wr_496  , wr_388  );
  nor  g846( wr_957  , wr_956  , wr_946  );
  nor  g847( wr_961  , wr_960  , G4088   );
  nor  g848( wr_1071 , wr_1070 , wr_1061 );
  nor  g849( wr_1074 , wr_1073 , G4089   );
  nor  g850( wr_1453 , wr_1452 , wr_1442 );
  nor  g851( wr_1457 , wr_1456 , G1689   );
  nor  g852( wr_1473 , wr_1472 , wr_1463 );
  nor  g853( wr_1476 , wr_1475 , G1691   );
  nor  g854( wr_1491 , wr_1490 , wr_946  );
  nor  g855( wr_1495 , wr_1494 , G4088   );
  nor  g856( wr_1510 , wr_1509 , wr_946  );
  nor  g857( wr_1514 , wr_1513 , G4088   );
  nor  g858( wr_1529 , wr_1528 , wr_946  );
  nor  g859( wr_1533 , wr_1532 , G4088   );
  nor  g860( wr_1548 , wr_1547 , wr_946  );
  nor  g861( wr_1552 , wr_1551 , G4088   );
  nor  g862( wr_1566 , wr_1565 , wr_1061 );
  nor  g863( wr_1569 , wr_1568 , G4089   );
  nor  g864( wr_1583 , wr_1582 , wr_1061 );
  nor  g865( wr_1586 , wr_1585 , G4089   );
  nor  g866( wr_1600 , wr_1599 , wr_1061 );
  nor  g867( wr_1603 , wr_1602 , G4089   );
  nor  g868( wr_1617 , wr_1616 , wr_1061 );
  nor  g869( wr_1620 , wr_1619 , G4089   );
  nor  g870( wr_1635 , wr_1634 , wr_1442 );
  nor  g871( wr_1639 , wr_1638 , G1689   );
  nor  g872( wr_1654 , wr_1653 , wr_1442 );
  nor  g873( wr_1658 , wr_1657 , G1689   );
  nor  g874( wr_1673 , wr_1672 , wr_1442 );
  nor  g875( wr_1677 , wr_1676 , G1689   );
  nor  g876( wr_1692 , wr_1691 , wr_1442 );
  nor  g877( wr_1696 , wr_1695 , G1689   );
  nor  g878( wr_1710 , wr_1709 , wr_1463 );
  nor  g879( wr_1713 , wr_1712 , G1691   );
  nor  g880( wr_1727 , wr_1726 , wr_1463 );
  nor  g881( wr_1730 , wr_1729 , G1691   );
  nor  g882( wr_1744 , wr_1743 , wr_1463 );
  nor  g883( wr_1747 , wr_1746 , G1691   );
  nor  g884( wr_1761 , wr_1760 , wr_1463 );
  nor  g885( wr_1764 , wr_1763 , G1691   );
  nor  g886( wr_1776 , wr_579  , wr_1775 );
  nor  g887( wr_1781 , wr_304  , G3717   );
  nor  g888( wr_1791 , wr_1790 , G3724   );
  nor  g889( wr_1861 , wr_1860 , wr_131  );
  nor  g890( wr_1928 , wr_1927 , wr_1061 );
  nor  g891( wr_1932 , wr_1931 , G4089   );
  nor  g892( wr_1946 , wr_1945 , wr_946  );
  nor  g893( wr_1949 , wr_1948 , G4088   );
  nor  g894( wr_1964 , wr_1963 , wr_946  );
  nor  g895( wr_1968 , wr_1967 , G4088   );
  nor  g896( wr_1983 , wr_1982 , wr_946  );
  nor  g897( wr_1987 , wr_1986 , G4088   );
  nor  g898( wr_2002 , wr_2001 , wr_946  );
  nor  g899( wr_2006 , wr_2005 , G4088   );
  nor  g900( wr_2020 , wr_2019 , wr_1061 );
  nor  g901( wr_2023 , wr_2022 , G4089   );
  nor  g902( wr_2037 , wr_2036 , wr_1061 );
  nor  g903( wr_2040 , wr_2039 , G4089   );
  nor  g904( wr_2054 , wr_2053 , wr_1061 );
  nor  g905( wr_2057 , wr_2056 , G4089   );
  nor  g906( wr_2072 , wr_2071 , wr_1442 );
  nor  g907( wr_2076 , wr_2075 , G1689   );
  nor  g908( wr_2091 , wr_2090 , wr_1442 );
  nor  g909( wr_2095 , wr_2094 , G1689   );
  nor  g910( wr_2110 , wr_2109 , wr_1442 );
  nor  g911( wr_2114 , wr_2113 , G1689   );
  nor  g912( wr_2129 , wr_2128 , wr_1442 );
  nor  g913( wr_2133 , wr_2132 , G1689   );
  nor  g914( wr_2147 , wr_2146 , wr_1463 );
  nor  g915( wr_2150 , wr_2149 , G1691   );
  nor  g916( wr_2164 , wr_2163 , wr_1463 );
  nor  g917( wr_2167 , wr_2166 , G1691   );
  nor  g918( wr_2181 , wr_2180 , wr_1463 );
  nor  g919( wr_2184 , wr_2183 , G1691   );
  nor  g920( wr_2198 , wr_2197 , wr_1463 );
  nor  g921( wr_2201 , wr_2200 , G1691   );
  nor  g922( wr_2475 , wr_2474 , G4091   );
  nor  g923( wr_2815 , wr_2814 , G4091   );
  nor  g924( wr_2846 , wr_2845 , wr_946  );
  nor  g925( wr_2850 , wr_2849 , G4088   );
  nor  g926( wr_2864 , wr_2863 , wr_1061 );
  nor  g927( wr_2867 , wr_2866 , G4089   );
  nor  g928( wr_157  , G809    , wr_156  );
  nor  g929( wr_170  , G809    , wr_169  );
  nor  g930( wr_181  , G809    , wr_180  );
  nor  g931( wr_192  , G809    , wr_191  );
  nor  g932( wr_137  , G809    , wr_134  );
  nor  g933( wr_144  , wr_143  , G809    );
  nor  g934( wr_150  , wr_149  , G809    );
  nor  g935( wr_155  , wr_154  , G809    );
  nor  g936( wr_483  , wr_482  , wr_452  );
  nor  g937( wr_491  , wr_490  , wr_404  );
  nor  g938( wr_507  , wr_506  , wr_436  );
  nor  g939( wr_521  , wr_520  , wr_318  );
  nor  g940( wr_529  , wr_528  , wr_334  );
  nor  g941( wr_537  , wr_536  , wr_366  );
  nor  g942( wr_553  , wr_552  , wr_350  );
  nor  g943( wr_569  , wr_568  , wr_285  );
  nor  g944( wr_586  , wr_585  , wr_267  );
  nor  g945( wr_603  , wr_602  , wr_601  );
  nor  g946( wr_608  , wr_607  , wr_202  );
  nor  g947( wr_615  , wr_614  , wr_218  );
  not  g948( wr_755  ,           wr_754  );
  not  g949( wr_782  ,           wr_781  );
  not  g950( wr_791  ,           wr_790  );
  not  g951( wr_808  ,           wr_807  );
  not  g952( wr_815  ,           wr_814  );
  not  g953( wr_842  ,           wr_841  );
  nor  g954( wr_1398 , wr_568  , G490    );
  nor  g955( wr_1312 , wr_490  , G422    );
  nor  g956( wr_2546 , wr_528  , G374    );
  not  g957( wr_762  ,           wr_761  );
  not  g958( wr_830  ,           wr_829  );
  nor  g959( wr_623  , wr_622  , wr_234  );
  not  g960( wr_777  ,           wr_776  );
  nor  g961( wr_545  , wr_544  , wr_420  );
  nor  g962( wr_499  , wr_498  , wr_388  );
  nor  g963( wr_2398 , wr_2397 , wr_2396 );
  nor  g964( wr_2411 , wr_2410 , wr_2409 );
  nor  g965( wr_2432 , wr_2431 , wr_2430 );
  nor  g966( wr_2404 , wr_2403 , wr_2400 );
  nor  g967( wr_2417 , wr_2416 , wr_2413 );
  nor  g968( wr_2438 , wr_2437 , wr_2434 );
  not  g969( wr_773  ,           wr_772  );
  nor  g970( wr_2717 , wr_2716 , wr_2715 );
  nor  g971( wr_2730 , wr_2729 , wr_2728 );
  nor  g972( wr_2747 , wr_2746 , wr_2745 );
  nor  g973( wr_2760 , wr_2759 , wr_2758 );
  nor  g974( wr_2723 , wr_2722 , wr_2719 );
  nor  g975( wr_2736 , wr_2735 , wr_2732 );
  nor  g976( wr_2753 , wr_2752 , wr_2749 );
  nor  g977( wr_2766 , wr_2765 , wr_2762 );
  nor  g978( wr_275  , wr_274  , wr_271  );
  nor  g979( wr_293  , wr_292  , wr_289  );
  nor  g980( wr_283  , wr_282  , wr_278  );
  nor  g981( wr_299  , wr_298  , wr_295  );
  nor  g982( wr_2777 , wr_2776 , wr_2775 );
  nor  g983( wr_396  , wr_395  , wr_392  );
  nor  g984( wr_2667 , wr_2666 , wr_2665 );
  nor  g985( wr_2680 , wr_2679 , wr_2678 );
  nor  g986( wr_2696 , wr_2695 , wr_2694 );
  nor  g987( wr_2783 , wr_2782 , wr_2779 );
  nor  g988( wr_402  , wr_401  , wr_398  );
  nor  g989( wr_2673 , wr_2672 , wr_2669 );
  nor  g990( wr_2686 , wr_2685 , wr_2682 );
  nor  g991( wr_2702 , wr_2701 , wr_2698 );
  nor  g992( wr_1254 , wr_506  , wr_480  );
  nor  g993( wr_1255 , wr_504  , wr_482  );
  nor  g994( wr_1263 , wr_1262 , wr_496  );
  nor  g995( wr_1264 , wr_1261 , wr_498  );
  nor  g996( wr_1267 , wr_542  , wr_490  );
  nor  g997( wr_1268 , wr_544  , wr_488  );
  nor  g998( wr_2386 , wr_1819 , wr_305  );
  nor  g999( wr_685  , wr_676  , G324    );
  nor g1000( wr_690  , wr_684  , wr_235  );
  nor g1001( wr_727  , wr_726  , wr_722  );
  nor g1002( wr_731  , wr_721  , wr_718  );
  nor g1003( wr_736  , wr_730  , wr_722  );
  not g1004( wr_682  ,           wr_681  );
  not g1005( wr_694  ,           wr_693  );
  not g1006( wr_740  ,           wr_739  );
  nor g1007( wr_210  , wr_209  , wr_206  );
  nor g1008( wr_226  , wr_225  , wr_222  );
  nor g1009( wr_242  , wr_241  , wr_238  );
  nor g1010( wr_216  , wr_215  , wr_212  );
  nor g1011( wr_232  , wr_231  , wr_228  );
  nor g1012( wr_248  , wr_247  , wr_244  );
  nor g1013( wr_1209 , wr_1208 , wr_597  );
  nor g1014( wr_1210 , wr_1207 , wr_598  );
  nor g1015( wr_1213 , wr_622  , wr_599  );
  nor g1016( wr_1217 , wr_614  , wr_606  );
  nor g1017( wr_1218 , wr_613  , wr_607  );
  nor g1018( wr_1243 , wr_526  , wr_520  );
  nor g1019( wr_1244 , wr_528  , wr_518  );
  nor g1020( wr_1246 , wr_552  , wr_534  );
  nor g1021( wr_1247 , wr_550  , wr_536  );
  nor g1022( wr_326  , wr_325  , wr_322  );
  nor g1023( wr_342  , wr_341  , wr_338  );
  nor g1024( wr_358  , wr_357  , wr_354  );
  nor g1025( wr_374  , wr_373  , wr_370  );
  nor g1026( wr_412  , wr_411  , wr_408  );
  nor g1027( wr_428  , wr_427  , wr_424  );
  nor g1028( wr_444  , wr_443  , wr_440  );
  nor g1029( wr_460  , wr_459  , wr_456  );
  nor g1030( wr_669  , wr_668  , wr_664  );
  nor g1031( wr_671  , wr_667  , wr_670  );
  nor g1032( wr_711  , wr_710  , wr_706  );
  nor g1033( wr_713  , wr_709  , wr_712  );
  nor g1034( wr_880  , wr_598  , G54     );
  nor g1035( wr_332  , wr_331  , wr_328  );
  nor g1036( wr_348  , wr_347  , wr_344  );
  nor g1037( wr_364  , wr_363  , wr_360  );
  nor g1038( wr_380  , wr_379  , wr_376  );
  nor g1039( wr_418  , wr_417  , wr_414  );
  nor g1040( wr_434  , wr_433  , wr_430  );
  nor g1041( wr_450  , wr_449  , wr_446  );
  nor g1042( wr_466  , wr_465  , wr_462  );
  nor g1043( wr_862  , wr_598  , G54     );
  nor g1044( wr_875  , wr_874  , G4092   );
  nor g1045( wr_1032 , wr_1031 , G4092   );
  nor g1046( wr_1820 , wr_1819 , G4092   );
  nor g1047( wr_806  , wr_580  , wr_575  );
  nor g1048( wr_1194 , wr_585  , wr_567  );
  nor g1049( wr_1195 , wr_584  , wr_568  );
  nor g1050( wr_1197 , wr_579  , wr_576  );
  not g1051( wr_1808 ,           wr_1807 );
  nor g1052( wr_310  , wr_309  , wr_305  );
  nor g1053( wr_634  , wr_580  , wr_576  );
  nor g1054( wr_1774 , wr_580  , G132    );
  nor g1055( wr_2887 , wr_2886 , wr_2882 );
  nor g1056( wr_2905 , wr_2904 , wr_2901 );
  not g1057( wr_162  ,           wr_161  );
  not g1058( wr_175  ,           wr_174  );
  not g1059( wr_186  ,           wr_185  );
  not g1060( wr_197  ,           wr_196  );
  not g1061( wr_751  ,           wr_750  );
  nor g1062( wr_962  , wr_961  , wr_957  );
  nor g1063( wr_1075 , wr_1074 , wr_1071 );
  nor g1064( wr_1458 , wr_1457 , wr_1453 );
  nor g1065( wr_1477 , wr_1476 , wr_1473 );
  nor g1066( wr_1496 , wr_1495 , wr_1491 );
  nor g1067( wr_1515 , wr_1514 , wr_1510 );
  nor g1068( wr_1534 , wr_1533 , wr_1529 );
  nor g1069( wr_1553 , wr_1552 , wr_1548 );
  nor g1070( wr_1570 , wr_1569 , wr_1566 );
  nor g1071( wr_1587 , wr_1586 , wr_1583 );
  nor g1072( wr_1604 , wr_1603 , wr_1600 );
  nor g1073( wr_1621 , wr_1620 , wr_1617 );
  nor g1074( wr_1640 , wr_1639 , wr_1635 );
  nor g1075( wr_1659 , wr_1658 , wr_1654 );
  nor g1076( wr_1678 , wr_1677 , wr_1673 );
  nor g1077( wr_1697 , wr_1696 , wr_1692 );
  nor g1078( wr_1714 , wr_1713 , wr_1710 );
  nor g1079( wr_1731 , wr_1730 , wr_1727 );
  nor g1080( wr_1748 , wr_1747 , wr_1744 );
  nor g1081( wr_1765 , wr_1764 , wr_1761 );
  not g1082( wr_1782 ,           wr_1781 );
  not g1083( wr_1862 ,           wr_1861 );
  nor g1084( wr_1933 , wr_1932 , wr_1928 );
  nor g1085( wr_1950 , wr_1949 , wr_1946 );
  nor g1086( wr_1969 , wr_1968 , wr_1964 );
  nor g1087( wr_1988 , wr_1987 , wr_1983 );
  nor g1088( wr_2007 , wr_2006 , wr_2002 );
  nor g1089( wr_2024 , wr_2023 , wr_2020 );
  nor g1090( wr_2041 , wr_2040 , wr_2037 );
  nor g1091( wr_2058 , wr_2057 , wr_2054 );
  nor g1092( wr_2077 , wr_2076 , wr_2072 );
  nor g1093( wr_2096 , wr_2095 , wr_2091 );
  nor g1094( wr_2115 , wr_2114 , wr_2110 );
  nor g1095( wr_2134 , wr_2133 , wr_2129 );
  nor g1096( wr_2151 , wr_2150 , wr_2147 );
  nor g1097( wr_2168 , wr_2167 , wr_2164 );
  nor g1098( wr_2185 , wr_2184 , wr_2181 );
  nor g1099( wr_2202 , wr_2201 , wr_2198 );
  nor g1100( wr_2476 , wr_2475 , wr_2471 );
  nor g1101( wr_2816 , wr_2815 , wr_2471 );
  nor g1102( wr_2851 , wr_2850 , wr_2846 );
  nor g1103( wr_2868 , wr_2867 , wr_2864 );
  not g1104( wr_158  ,           wr_157  );
  not g1105( wr_171  ,           wr_170  );
  not g1106( wr_182  ,           wr_181  );
  not g1107( wr_193  ,           wr_192  );
  not g1108( G656    ,           wr_137  );
  not g1109( G636    ,           wr_144  );
  not g1110( G704    ,           wr_150  );
  not g1111( G820    ,           wr_155  );
  not g1112( G717    ,           wr_150  );
  nor g1113( wr_484  , wr_483  , wr_481  );
  nor g1114( wr_492  , wr_491  , wr_489  );
  nor g1115( wr_508  , wr_507  , wr_505  );
  nor g1116( wr_522  , wr_521  , wr_519  );
  nor g1117( wr_530  , wr_529  , wr_527  );
  nor g1118( wr_538  , wr_537  , wr_535  );
  nor g1119( wr_554  , wr_553  , wr_551  );
  nor g1120( wr_571  , wr_570  , wr_569  );
  nor g1121( wr_588  , wr_587  , wr_586  );
  nor g1122( wr_610  , wr_609  , wr_608  );
  nor g1123( wr_617  , wr_616  , wr_615  );
  nor g1124( wr_834  , wr_603  , wr_597  );
  not g1125( wr_1400 ,           wr_1398 );
  nor g1126( wr_816  , wr_815  , wr_576  );
  not g1127( wr_1314 ,           wr_1312 );
  not g1128( wr_2549 ,           wr_2546 );
  nor g1129( wr_831  , wr_830  , wr_603  );
  nor g1130( wr_625  , wr_624  , wr_623  );
  nor g1131( wr_843  , wr_842  , wr_603  );
  nor g1132( wr_546  , wr_545  , wr_543  );
  nor g1133( wr_500  , wr_499  , wr_497  );
  nor g1134( wr_809  , wr_808  , wr_576  );
  not g1135( wr_2399 ,           wr_2398 );
  not g1136( wr_2412 ,           wr_2411 );
  not g1137( wr_2433 ,           wr_2432 );
  not g1138( wr_2718 ,           wr_2717 );
  not g1139( wr_2731 ,           wr_2730 );
  not g1140( wr_2748 ,           wr_2747 );
  not g1141( wr_2761 ,           wr_2760 );
  not g1142( wr_276  ,           wr_275  );
  not g1143( wr_294  ,           wr_293  );
  not g1144( wr_1021 ,           wr_603  );
  not g1145( wr_2778 ,           wr_2777 );
  not g1146( wr_397  ,           wr_396  );
  not g1147( wr_2668 ,           wr_2667 );
  not g1148( wr_2681 ,           wr_2680 );
  not g1149( wr_2697 ,           wr_2696 );
  nor g1150( wr_1256 , wr_1255 , wr_1254 );
  nor g1151( wr_1265 , wr_1264 , wr_1263 );
  nor g1152( wr_1269 , wr_1268 , wr_1267 );
  nor g1153( wr_2388 , wr_2387 , wr_2386 );
  not g1154( wr_686  ,           wr_685  );
  not g1155( wr_691  ,           wr_690  );
  not g1156( wr_728  ,           wr_727  );
  not g1157( wr_732  ,           wr_731  );
  not g1158( wr_737  ,           wr_736  );
  nor g1159( wr_683  , wr_682  , wr_676  );
  nor g1160( wr_695  , wr_694  , wr_680  );
  nor g1161( wr_741  , wr_740  , wr_726  );
  not g1162( wr_211  ,           wr_210  );
  not g1163( wr_227  ,           wr_226  );
  not g1164( wr_243  ,           wr_242  );
  nor g1165( wr_1211 , wr_1210 , wr_1209 );
  nor g1166( wr_1215 , wr_1214 , wr_1213 );
  nor g1167( wr_1219 , wr_1218 , wr_1217 );
  nor g1168( wr_1245 , wr_1244 , wr_1243 );
  nor g1169( wr_1248 , wr_1247 , wr_1246 );
  not g1170( wr_327  ,           wr_326  );
  not g1171( wr_343  ,           wr_342  );
  not g1172( wr_359  ,           wr_358  );
  not g1173( wr_375  ,           wr_374  );
  not g1174( wr_413  ,           wr_412  );
  not g1175( wr_429  ,           wr_428  );
  not g1176( wr_445  ,           wr_444  );
  not g1177( wr_461  ,           wr_460  );
  nor g1178( wr_672  , wr_671  , wr_669  );
  nor g1179( wr_714  , wr_713  , wr_711  );
  not g1180( wr_881  ,           wr_880  );
  nor g1181( wr_865  , wr_864  , wr_862  );
  not g1182( wr_876  ,           wr_875  );
  not g1183( wr_1033 ,           wr_1032 );
  not g1184( wr_1821 ,           wr_1820 );
  nor g1185( wr_1196 , wr_1195 , wr_1194 );
  nor g1186( wr_1198 , wr_1197 , wr_806  );
  nor g1187( wr_1809 , wr_1808 , G4091   );
  not g1188( wr_311  ,           wr_310  );
  not g1189( wr_635  ,           wr_634  );
  nor g1190( wr_1777 , wr_1776 , wr_1774 );
  not g1191( wr_2888 ,           wr_2887 );
  not g1192( wr_2906 ,           wr_2905 );
  nor g1193( wr_163  , wr_162  , G2358   );
  nor g1194( wr_176  , wr_175  , G2358   );
  nor g1195( wr_187  , wr_186  , G2358   );
  nor g1196( wr_198  , wr_197  , G2358   );
  not g1197( wr_963  ,           wr_962  );
  not g1198( wr_1076 ,           wr_1075 );
  not g1199( wr_1459 ,           wr_1458 );
  not g1200( wr_1478 ,           wr_1477 );
  not g1201( wr_1497 ,           wr_1496 );
  not g1202( wr_1516 ,           wr_1515 );
  not g1203( wr_1535 ,           wr_1534 );
  not g1204( wr_1554 ,           wr_1553 );
  not g1205( wr_1571 ,           wr_1570 );
  not g1206( wr_1588 ,           wr_1587 );
  not g1207( wr_1605 ,           wr_1604 );
  not g1208( wr_1622 ,           wr_1621 );
  not g1209( wr_1641 ,           wr_1640 );
  not g1210( wr_1660 ,           wr_1659 );
  not g1211( wr_1679 ,           wr_1678 );
  not g1212( wr_1698 ,           wr_1697 );
  not g1213( wr_1715 ,           wr_1714 );
  not g1214( wr_1732 ,           wr_1731 );
  not g1215( wr_1749 ,           wr_1748 );
  not g1216( wr_1766 ,           wr_1765 );
  nor g1217( wr_1783 , wr_1782 , G3724   );
  nor g1218( wr_1863 , wr_1862 , G851    );
  not g1219( wr_1934 ,           wr_1933 );
  not g1220( wr_1951 ,           wr_1950 );
  not g1221( wr_1970 ,           wr_1969 );
  not g1222( wr_1989 ,           wr_1988 );
  not g1223( wr_2008 ,           wr_2007 );
  not g1224( wr_2025 ,           wr_2024 );
  not g1225( wr_2042 ,           wr_2041 );
  not g1226( wr_2059 ,           wr_2058 );
  not g1227( wr_2078 ,           wr_2077 );
  not g1228( wr_2097 ,           wr_2096 );
  not g1229( wr_2116 ,           wr_2115 );
  not g1230( wr_2135 ,           wr_2134 );
  not g1231( wr_2152 ,           wr_2151 );
  not g1232( wr_2169 ,           wr_2168 );
  not g1233( wr_2186 ,           wr_2185 );
  not g1234( wr_2203 ,           wr_2202 );
  not g1235( wr_2477 ,           wr_2476 );
  not g1236( wr_2817 ,           wr_2816 );
  not g1237( wr_2852 ,           wr_2851 );
  not g1238( wr_2869 ,           wr_2868 );
  nor g1239( wr_159  , wr_158  , wr_139  );
  nor g1240( wr_172  , wr_171  , wr_139  );
  nor g1241( wr_183  , wr_182  , wr_139  );
  nor g1242( wr_194  , wr_193  , wr_139  );
  nor g1243( wr_783  , wr_782  , wr_554  );
  not g1244( wr_835  ,           wr_834  );
  nor g1245( wr_930  , wr_576  , wr_571  );
  nor g1246( wr_933  , wr_588  , wr_576  );
  nor g1247( wr_967  , wr_610  , wr_603  );
  nor g1248( wr_970  , wr_617  , wr_603  );
  nor g1249( wr_1005 , wr_842  , wr_610  );
  nor g1250( wr_1011 , wr_617  , wr_597  );
  nor g1251( wr_1080 , wr_554  , wr_538  );
  nor g1252( wr_1083 , wr_554  , wr_522  );
  nor g1253( wr_1118 , wr_791  , wr_538  );
  nor g1254( wr_1124 , wr_782  , wr_522  );
  nor g1255( wr_1331 , wr_508  , wr_492  );
  nor g1256( wr_1334 , wr_508  , wr_484  );
  nor g1257( wr_1349 , wr_755  , wr_484  );
  nor g1258( wr_1358 , wr_492  , wr_484  );
  nor g1259( wr_1408 , wr_808  , wr_588  );
  nor g1260( wr_1416 , wr_588  , wr_571  );
  nor g1261( wr_2263 , wr_617  , wr_598  );
  nor g1262( wr_2537 , wr_530  , wr_522  );
  nor g1263( wr_763  , wr_762  , wr_508  );
  nor g1264( wr_778  , wr_777  , wr_554  );
  not g1265( wr_844  ,           wr_843  );
  not g1266( wr_1389 ,           wr_571  );
  nor g1267( wr_792  , wr_791  , wr_554  );
  not g1268( wr_1303 ,           wr_492  );
  not g1269( wr_1394 ,           wr_588  );
  not g1270( wr_832  ,           wr_831  );
  not g1271( wr_901  ,           wr_530  );
  nor g1272( wr_640  , wr_625  , wr_603  );
  not g1273( wr_883  ,           wr_617  );
  not g1274( wr_1308 ,           wr_484  );
  nor g1275( wr_555  , wr_554  , wr_546  );
  nor g1276( wr_626  , wr_625  , wr_617  );
  nor g1277( wr_654  , wr_546  , wr_522  );
  not g1278( wr_1178 ,           wr_522  );
  nor g1279( wr_756  , wr_755  , wr_508  );
  not g1280( wr_989  ,           wr_625  );
  not g1281( wr_1325 ,           wr_500  );
  not g1282( wr_810  ,           wr_809  );
  nor g1283( wr_827  , wr_826  , wr_625  );
  not g1284( wr_1102 ,           wr_546  );
  nor g1285( wr_2405 , wr_2404 , wr_2399 );
  nor g1286( wr_2418 , wr_2417 , wr_2412 );
  nor g1287( wr_2439 , wr_2438 , wr_2433 );
  nor g1288( wr_774  , wr_773  , wr_546  );
  not g1289( wr_1045 ,           wr_610  );
  not g1290( wr_1352 ,           wr_508  );
  nor g1291( wr_1006 , wr_617  , wr_610  );
  nor g1292( wr_2724 , wr_2723 , wr_2718 );
  nor g1293( wr_2737 , wr_2736 , wr_2731 );
  nor g1294( wr_2754 , wr_2753 , wr_2748 );
  nor g1295( wr_2767 , wr_2766 , wr_2761 );
  not g1296( wr_1158 ,           wr_538  );
  nor g1297( wr_284  , wr_283  , wr_276  );
  nor g1298( wr_300  , wr_299  , wr_294  );
  nor g1299( wr_1119 , wr_538  , wr_522  );
  nor g1300( wr_2784 , wr_2783 , wr_2778 );
  nor g1301( wr_403  , wr_402  , wr_397  );
  nor g1302( wr_1037 , wr_617  , wr_863  );
  not g1303( wr_1134 ,           wr_554  );
  nor g1304( wr_2674 , wr_2673 , wr_2668 );
  nor g1305( wr_2687 , wr_2686 , wr_2681 );
  nor g1306( wr_2703 , wr_2702 , wr_2697 );
  nor g1307( wr_1313 , wr_1312 , wr_484  );
  nor g1308( wr_1399 , wr_1398 , wr_588  );
  nor g1309( wr_1150 , wr_522  , wr_900  );
  not g1310( wr_1257 ,           wr_1256 );
  not g1311( wr_1266 ,           wr_1265 );
  not g1312( wr_1273 ,           wr_1269 );
  nor g1313( wr_1307 , wr_754  , wr_484  );
  nor g1314( wr_1393 , wr_807  , wr_588  );
  not g1315( wr_2389 ,           wr_2388 );
  nor g1316( wr_687  , wr_686  , wr_684  );
  nor g1317( wr_692  , wr_691  , wr_675  );
  nor g1318( wr_729  , wr_728  , wr_718  );
  nor g1319( wr_733  , wr_732  , wr_730  );
  nor g1320( wr_738  , wr_737  , wr_717  );
  nor g1321( wr_1282 , wr_1265 , wr_1256 );
  nor g1322( wr_217  , wr_216  , wr_211  );
  nor g1323( wr_233  , wr_232  , wr_227  );
  nor g1324( wr_249  , wr_248  , wr_243  );
  nor g1325( wr_1174 , wr_530  , wr_900  );
  not g1326( wr_1212 ,           wr_1211 );
  not g1327( wr_1216 ,           wr_1215 );
  not g1328( wr_1223 ,           wr_1219 );
  not g1329( wr_1249 ,           wr_1248 );
  not g1330( wr_1251 ,           wr_1245 );
  nor g1331( wr_333  , wr_332  , wr_327  );
  nor g1332( wr_349  , wr_348  , wr_343  );
  nor g1333( wr_365  , wr_364  , wr_359  );
  nor g1334( wr_381  , wr_380  , wr_375  );
  nor g1335( wr_419  , wr_418  , wr_413  );
  nor g1336( wr_435  , wr_434  , wr_429  );
  nor g1337( wr_451  , wr_450  , wr_445  );
  nor g1338( wr_467  , wr_466  , wr_461  );
  not g1339( wr_701  ,           wr_672  );
  not g1340( wr_747  ,           wr_714  );
  nor g1341( wr_882  , wr_881  , wr_617  );
  nor g1342( wr_1232 , wr_1215 , wr_1211 );
  nor g1343( wr_866  , wr_865  , G4092   );
  nor g1344( wr_877  , wr_876  , G4091   );
  nor g1345( wr_899  , wr_530  , G4      );
  nor g1346( wr_1034 , wr_1033 , G4091   );
  nor g1347( wr_1822 , wr_1821 , G4091   );
  not g1348( wr_817  ,           wr_816  );
  not g1349( wr_1199 ,           wr_1198 );
  not g1350( wr_1201 ,           wr_1196 );
  nor g1351( wr_1810 , wr_1809 , wr_1806 );
  nor g1352( wr_509  , wr_508  , wr_500  );
  nor g1353( wr_589  , wr_588  , wr_580  );
  nor g1354( wr_648  , wr_500  , wr_484  );
  nor g1355( wr_636  , wr_635  , wr_571  );
  nor g1356( wr_752  , wr_751  , wr_500  );
  nor g1357( wr_1778 , wr_1777 , G3717   );
  nor g1358( wr_166  , wr_165  , wr_163  );
  nor g1359( wr_177  , wr_176  , wr_165  );
  nor g1360( wr_188  , wr_187  , wr_165  );
  nor g1361( wr_199  , wr_198  , wr_165  );
  not g1362( wr_1384 ,           wr_865  );
  not g1363( wr_1798 ,           wr_1777 );
  not g1364( wr_1864 ,           wr_1863 );
  not g1365( wr_784  ,           wr_783  );
  not g1366( wr_931  ,           wr_930  );
  not g1367( wr_934  ,           wr_933  );
  not g1368( wr_968  ,           wr_967  );
  not g1369( wr_971  ,           wr_970  );
  nor g1370( wr_977  , wr_835  , wr_617  );
  not g1371( wr_1012 ,           wr_1011 );
  not g1372( wr_1081 ,           wr_1080 );
  not g1373( wr_1084 ,           wr_1083 );
  not g1374( wr_1125 ,           wr_1124 );
  not g1375( wr_1332 ,           wr_1331 );
  not g1376( wr_1335 ,           wr_1334 );
  nor g1377( wr_1350 , wr_1349 , wr_761  );
  nor g1378( wr_1409 , wr_1408 , wr_814  );
  nor g1379( wr_2213 , wr_1011 , wr_841  );
  not g1380( wr_2265 ,           wr_2263 );
  not g1381( wr_2539 ,           wr_2537 );
  nor g1382( wr_2487 , wr_1124 , wr_790  );
  nor g1383( wr_836  , wr_835  , wr_625  );
  nor g1384( wr_845  , wr_844  , wr_610  );
  not g1385( wr_793  ,           wr_792  );
  nor g1386( wr_833  , wr_832  , wr_625  );
  not g1387( wr_641  ,           wr_640  );
  not g1388( wr_779  ,           wr_778  );
  not g1389( wr_556  ,           wr_555  );
  not g1390( wr_627  ,           wr_626  );
  not g1391( wr_655  ,           wr_654  );
  not g1392( wr_757  ,           wr_756  );
  nor g1393( wr_811  , wr_810  , wr_588  );
  not g1394( wr_2406 ,           wr_2405 );
  not g1395( wr_2420 ,           wr_2418 );
  not g1396( wr_2441 ,           wr_2439 );
  nor g1397( wr_1359 , wr_1358 , wr_761  );
  nor g1398( wr_1417 , wr_1416 , wr_814  );
  nor g1399( wr_2440 , wr_2439 , wr_2427 );
  not g1400( wr_1007 ,           wr_1006 );
  not g1401( wr_2725 ,           wr_2724 );
  not g1402( wr_2739 ,           wr_2737 );
  not g1403( wr_2755 ,           wr_2754 );
  not g1404( wr_2769 ,           wr_2767 );
  not g1405( wr_1120 ,           wr_1119 );
  not g1406( wr_1832 ,           wr_284  );
  not g1407( wr_1845 ,           wr_300  );
  not g1408( wr_2788 ,           wr_2784 );
  not g1409( wr_1038 ,           wr_1037 );
  nor g1410( wr_1315 , wr_1314 , wr_1308 );
  nor g1411( wr_1401 , wr_1400 , wr_1394 );
  not g1412( wr_1874 ,           wr_403  );
  not g1413( wr_2675 ,           wr_2674 );
  not g1414( wr_2689 ,           wr_2687 );
  not g1415( wr_2704 ,           wr_2703 );
  nor g1416( wr_1309 , wr_755  , wr_1308 );
  nor g1417( wr_1395 , wr_808  , wr_1394 );
  not g1418( wr_1151 ,           wr_1150 );
  nor g1419( wr_1270 , wr_1269 , wr_1266 );
  nor g1420( wr_1274 , wr_1265 , wr_1257 );
  nor g1421( wr_1279 , wr_1273 , wr_1266 );
  nor g1422( wr_688  , wr_687  , wr_683  );
  nor g1423( wr_696  , wr_695  , wr_692  );
  nor g1424( wr_734  , wr_733  , wr_729  );
  nor g1425( wr_742  , wr_741  , wr_738  );
  not g1426( wr_1283 ,           wr_1282 );
  not g1427( wr_893  ,           wr_233  );
  not g1428( wr_999  ,           wr_249  );
  not g1429( wr_1055 ,           wr_217  );
  nor g1430( wr_884  , wr_880  , wr_883  );
  nor g1431( wr_1175 , wr_1174 , wr_781  );
  nor g1432( wr_1220 , wr_1219 , wr_1216 );
  nor g1433( wr_1224 , wr_1215 , wr_1212 );
  nor g1434( wr_1229 , wr_1223 , wr_1216 );
  nor g1435( wr_1250 , wr_1249 , wr_1245 );
  nor g1436( wr_1252 , wr_1248 , wr_1251 );
  not g1437( wr_911  ,           wr_349  );
  not g1438( wr_1112 ,           wr_435  );
  not g1439( wr_1144 ,           wr_365  );
  not g1440( wr_1168 ,           wr_381  );
  not g1441( wr_1188 ,           wr_333  );
  not g1442( wr_1233 ,           wr_1232 );
  not g1443( wr_1887 ,           wr_451  );
  not g1444( wr_1900 ,           wr_467  );
  not g1445( wr_1913 ,           wr_419  );
  nor g1446( wr_902  , wr_901  , wr_900  );
  not g1447( wr_764  ,           wr_763  );
  not g1448( wr_867  ,           wr_866  );
  nor g1449( wr_878  , wr_877  , wr_873  );
  nor g1450( wr_1035 , wr_1034 , wr_1030 );
  nor g1451( wr_1823 , wr_1822 , wr_1818 );
  nor g1452( wr_468  , wr_467  , wr_451  );
  nor g1453( wr_818  , wr_817  , wr_580  );
  nor g1454( wr_1200 , wr_1199 , wr_1196 );
  nor g1455( wr_1202 , wr_1198 , wr_1201 );
  not g1456( wr_1811 ,           wr_1810 );
  not g1457( wr_510  ,           wr_509  );
  not g1458( wr_590  ,           wr_589  );
  not g1459( wr_649  ,           wr_648  );
  nor g1460( wr_255  , wr_254  , wr_249  );
  nor g1461( wr_312  , wr_311  , wr_300  );
  nor g1462( wr_382  , wr_381  , wr_365  );
  not g1463( wr_637  ,           wr_636  );
  not g1464( wr_1779 ,           wr_1778 );
  not g1465( wr_167  ,           wr_166  );
  not g1466( wr_178  ,           wr_177  );
  not g1467( wr_189  ,           wr_188  );
  not g1468( wr_200  ,           wr_199  );
  nor g1469( wr_1865 , wr_1864 , G848    );
  nor g1470( wr_932  , wr_931  , wr_588  );
  nor g1471( wr_935  , wr_934  , wr_808  );
  nor g1472( wr_969  , wr_968  , wr_842  );
  not g1473( wr_978  ,           wr_977  );
  nor g1474( wr_1013 , wr_1012 , wr_610  );
  nor g1475( wr_1090 , wr_784  , wr_522  );
  nor g1476( wr_1126 , wr_1125 , wr_538  );
  nor g1477( wr_1333 , wr_1332 , wr_484  );
  nor g1478( wr_1336 , wr_1335 , wr_755  );
  not g1479( wr_1353 ,           wr_1350 );
  not g1480( wr_1411 ,           wr_1409 );
  nor g1481( wr_2253 , wr_971  , wr_598  );
  nor g1482( wr_2266 , wr_2265 , wr_610  );
  nor g1483( wr_2527 , wr_1084 , wr_530  );
  nor g1484( wr_2540 , wr_2539 , wr_538  );
  nor g1485( wr_1082 , wr_1081 , wr_791  );
  not g1486( wr_2214 ,           wr_2213 );
  nor g1487( wr_2337 , wr_1409 , wr_808  );
  not g1488( wr_2488 ,           wr_2487 );
  nor g1489( wr_2617 , wr_1350 , wr_755  );
  not g1490( wr_837  ,           wr_836  );
  nor g1491( wr_785  , wr_784  , wr_546  );
  not g1492( wr_846  ,           wr_845  );
  nor g1493( wr_794  , wr_793  , wr_538  );
  nor g1494( wr_642  , wr_641  , wr_610  );
  nor g1495( wr_780  , wr_779  , wr_546  );
  nor g1496( wr_557  , wr_556  , wr_538  );
  nor g1497( wr_628  , wr_627  , wr_610  );
  nor g1498( wr_656  , wr_655  , wr_538  );
  nor g1499( wr_758  , wr_757  , wr_484  );
  nor g1500( wr_972  , wr_971  , wr_610  );
  nor g1501( wr_917  , wr_811  , wr_576  );
  nor g1502( wr_1085 , wr_1084 , wr_538  );
  nor g1503( wr_2419 , wr_2418 , wr_2406 );
  nor g1504( wr_2421 , wr_2420 , wr_2405 );
  nor g1505( wr_2442 , wr_2441 , wr_2426 );
  not g1506( wr_1360 ,           wr_1359 );
  not g1507( wr_1418 ,           wr_1417 );
  nor g1508( wr_1008 , wr_1007 , wr_863  );
  nor g1509( wr_2738 , wr_2737 , wr_2725 );
  nor g1510( wr_2740 , wr_2739 , wr_2724 );
  nor g1511( wr_2768 , wr_2767 , wr_2755 );
  nor g1512( wr_2770 , wr_2769 , wr_2754 );
  nor g1513( wr_1351 , wr_1350 , wr_508  );
  nor g1514( wr_1410 , wr_1409 , wr_576  );
  nor g1515( wr_1121 , wr_1120 , wr_900  );
  nor g1516( wr_2383 , wr_1845 , wr_284  );
  nor g1517( wr_2384 , wr_300  , wr_1832 );
  nor g1518( wr_1039 , wr_1038 , wr_598  );
  nor g1519( wr_1316 , wr_1315 , wr_1313 );
  nor g1520( wr_1402 , wr_1401 , wr_1399 );
  nor g1521( wr_2688 , wr_2687 , wr_2675 );
  nor g1522( wr_2690 , wr_2689 , wr_2674 );
  nor g1523( wr_2705 , wr_2704 , wr_403  );
  nor g1524( wr_2706 , wr_2703 , wr_1874 );
  nor g1525( wr_1310 , wr_1309 , wr_1307 );
  nor g1526( wr_1396 , wr_1395 , wr_1393 );
  nor g1527( wr_1152 , wr_1151 , wr_530  );
  not g1528( wr_1271 ,           wr_1270 );
  not g1529( wr_1275 ,           wr_1274 );
  not g1530( wr_1280 ,           wr_1279 );
  not g1531( wr_689  ,           wr_688  );
  not g1532( wr_697  ,           wr_696  );
  not g1533( wr_735  ,           wr_734  );
  not g1534( wr_743  ,           wr_742  );
  nor g1535( wr_1284 , wr_1283 , wr_1269 );
  nor g1536( wr_894  , wr_893  , G4092   );
  nor g1537( wr_1000 , wr_999  , G4092   );
  nor g1538( wr_1056 , wr_1055 , G4092   );
  nor g1539( wr_1833 , wr_1832 , G4092   );
  nor g1540( wr_1846 , wr_1845 , G4092   );
  nor g1541( wr_885  , wr_884  , wr_882  );
  not g1542( wr_1176 ,           wr_1175 );
  not g1543( wr_1221 ,           wr_1220 );
  not g1544( wr_1225 ,           wr_1224 );
  not g1545( wr_1230 ,           wr_1229 );
  nor g1546( wr_1253 , wr_1252 , wr_1250 );
  nor g1547( wr_912  , wr_911  , G4092   );
  nor g1548( wr_1113 , wr_1112 , G4092   );
  nor g1549( wr_1145 , wr_1144 , G4092   );
  nor g1550( wr_1169 , wr_1168 , G4092   );
  nor g1551( wr_1179 , wr_1175 , wr_1178 );
  nor g1552( wr_1189 , wr_1188 , G4092   );
  nor g1553( wr_1234 , wr_1233 , wr_1219 );
  nor g1554( wr_1875 , wr_1874 , G4092   );
  nor g1555( wr_1888 , wr_1887 , G4092   );
  nor g1556( wr_1901 , wr_1900 , G4092   );
  nor g1557( wr_1914 , wr_1913 , G4092   );
  not g1558( wr_812  ,           wr_811  );
  nor g1559( wr_903  , wr_902  , wr_899  );
  nor g1560( wr_765  , wr_764  , wr_500  );
  nor g1561( wr_868  , wr_867  , wr_861  );
  not g1562( wr_879  ,           wr_878  );
  not g1563( wr_1036 ,           wr_1035 );
  not g1564( wr_1824 ,           wr_1823 );
  not g1565( wr_469  ,           wr_468  );
  nor g1566( wr_1203 , wr_1202 , wr_1200 );
  nor g1567( wr_511  , wr_510  , wr_492  );
  nor g1568( wr_591  , wr_590  , wr_576  );
  nor g1569( wr_650  , wr_649  , wr_508  );
  not g1570( wr_256  ,           wr_255  );
  not g1571( wr_313  ,           wr_312  );
  not g1572( wr_383  ,           wr_382  );
  nor g1573( wr_638  , wr_637  , wr_588  );
  nor g1574( wr_1780 , wr_1779 , wr_1773 );
  nor g1575( wr_168  , wr_167  , wr_159  );
  nor g1576( wr_179  , wr_178  , wr_172  );
  nor g1577( wr_190  , wr_189  , wr_183  );
  nor g1578( wr_201  , wr_200  , wr_194  );
  not g1579( wr_1866 ,           wr_1865 );
  nor g1580( wr_936  , wr_935  , wr_932  );
  nor g1581( wr_979  , wr_978  , wr_610  );
  not g1582( wr_1091 ,           wr_1090 );
  nor g1583( wr_1337 , wr_1336 , wr_1333 );
  nor g1584( wr_2215 , wr_1013 , wr_829  );
  not g1585( wr_2254 ,           wr_2253 );
  nor g1586( wr_2267 , wr_2266 , wr_1013 );
  nor g1587( wr_2304 , wr_1416 , wr_1411 );
  nor g1588( wr_2332 , wr_935  , wr_576  );
  nor g1589( wr_2489 , wr_1126 , wr_776  );
  not g1590( wr_2528 ,           wr_2527 );
  nor g1591( wr_2541 , wr_2540 , wr_1126 );
  nor g1592( wr_2336 , wr_1411 , wr_807  );
  nor g1593( wr_2584 , wr_1358 , wr_1353 );
  nor g1594( wr_2264 , wr_2263 , wr_2214 );
  nor g1595( wr_2612 , wr_1336 , wr_750  );
  nor g1596( wr_2616 , wr_1353 , wr_754  );
  nor g1597( wr_2538 , wr_2537 , wr_2488 );
  nor g1598( wr_838  , wr_837  , wr_617  );
  not g1599( wr_786  ,           wr_785  );
  nor g1600( wr_847  , wr_846  , wr_625  );
  not g1601( wr_795  ,           wr_794  );
  not g1602( wr_643  ,           wr_642  );
  not g1603( wr_558  ,           wr_557  );
  not g1604( wr_629  ,           wr_628  );
  not g1605( wr_657  ,           wr_656  );
  not g1606( wr_973  ,           wr_972  );
  nor g1607( wr_1321 , wr_758  , wr_750  );
  not g1608( wr_918  ,           wr_917  );
  not g1609( wr_1086 ,           wr_1085 );
  nor g1610( wr_2422 , wr_2421 , wr_2419 );
  nor g1611( wr_2443 , wr_2442 , wr_2440 );
  nor g1612( wr_1361 , wr_1360 , wr_1349 );
  nor g1613( wr_1419 , wr_1418 , wr_1408 );
  not g1614( wr_1009 ,           wr_1008 );
  nor g1615( wr_1354 , wr_1353 , wr_1352 );
  nor g1616( wr_1412 , wr_1411 , wr_575  );
  nor g1617( wr_2741 , wr_2740 , wr_2738 );
  nor g1618( wr_2771 , wr_2770 , wr_2768 );
  not g1619( wr_1122 ,           wr_1121 );
  nor g1620( wr_2385 , wr_2384 , wr_2383 );
  nor g1621( wr_1040 , wr_1039 , wr_841  );
  not g1622( wr_1317 ,           wr_1316 );
  not g1623( wr_1403 ,           wr_1402 );
  nor g1624( wr_2691 , wr_2690 , wr_2688 );
  nor g1625( wr_2707 , wr_2706 , wr_2705 );
  nor g1626( wr_1153 , wr_1152 , wr_790  );
  nor g1627( wr_1272 , wr_1271 , wr_1257 );
  nor g1628( wr_1276 , wr_1275 , wr_1273 );
  nor g1629( wr_1281 , wr_1280 , wr_1256 );
  nor g1630( wr_698  , wr_697  , wr_689  );
  nor g1631( wr_744  , wr_743  , wr_735  );
  not g1632( wr_895  ,           wr_894  );
  not g1633( wr_1001 ,           wr_1000 );
  not g1634( wr_1057 ,           wr_1056 );
  not g1635( wr_1834 ,           wr_1833 );
  not g1636( wr_1847 ,           wr_1846 );
  nor g1637( wr_886  , wr_885  , G4092   );
  nor g1638( wr_1177 , wr_1176 , wr_522  );
  nor g1639( wr_1222 , wr_1221 , wr_1212 );
  nor g1640( wr_1226 , wr_1225 , wr_1223 );
  nor g1641( wr_1231 , wr_1230 , wr_1211 );
  not g1642( wr_1290 ,           wr_1253 );
  not g1643( wr_759  ,           wr_758  );
  not g1644( wr_913  ,           wr_912  );
  not g1645( wr_1114 ,           wr_1113 );
  not g1646( wr_1146 ,           wr_1145 );
  not g1647( wr_1170 ,           wr_1169 );
  not g1648( wr_1190 ,           wr_1189 );
  not g1649( wr_1876 ,           wr_1875 );
  not g1650( wr_1889 ,           wr_1888 );
  not g1651( wr_1902 ,           wr_1901 );
  not g1652( wr_1915 ,           wr_1914 );
  nor g1653( wr_813  , wr_812  , wr_580  );
  nor g1654( wr_904  , wr_903  , G4092   );
  nor g1655( G822    , wr_879  , wr_868  );
  nor g1656( wr_470  , wr_469  , wr_435  );
  not g1657( wr_1240 ,           wr_1203 );
  not g1658( wr_512  ,           wr_511  );
  not g1659( wr_592  ,           wr_591  );
  not g1660( wr_651  ,           wr_650  );
  nor g1661( wr_257  , wr_256  , wr_233  );
  nor g1662( wr_314  , wr_313  , wr_284  );
  nor g1663( wr_384  , wr_383  , wr_349  );
  not g1664( wr_639  ,           wr_638  );
  not g1665( wr_1294 ,           wr_903  );
  not g1666( wr_1383 ,           wr_885  );
  nor g1667( G639    , wr_168  , wr_124  );
  nor g1668( G673    , wr_179  , wr_124  );
  nor g1669( G707    , wr_190  , wr_124  );
  nor g1670( G715    , wr_201  , wr_124  );
  not g1671( wr_937  ,           wr_936  );
  nor g1672( wr_1092 , wr_1091 , wr_538  );
  nor g1673( wr_2207 , wr_979  , wr_969  );
  not g1674( wr_2216 ,           wr_2215 );
  nor g1675( wr_2255 , wr_2254 , wr_610  );
  not g1676( wr_2268 ,           wr_2267 );
  not g1677( wr_2306 ,           wr_2304 );
  not g1678( wr_2490 ,           wr_2489 );
  nor g1679( wr_2529 , wr_2528 , wr_538  );
  not g1680( wr_2542 ,           wr_2541 );
  not g1681( wr_1338 ,           wr_1337 );
  nor g1682( wr_2305 , wr_2304 , wr_1398 );
  not g1683( wr_2333 ,           wr_2332 );
  nor g1684( wr_2338 , wr_2337 , wr_2336 );
  not g1685( wr_2586 ,           wr_2584 );
  not g1686( wr_2274 ,           wr_2264 );
  nor g1687( wr_2585 , wr_2584 , wr_1312 );
  not g1688( wr_2613 ,           wr_2612 );
  nor g1689( wr_2618 , wr_2617 , wr_2616 );
  not g1690( wr_2554 ,           wr_2538 );
  not g1691( wr_839  ,           wr_838  );
  nor g1692( wr_787  , wr_786  , wr_522  );
  nor g1693( wr_796  , wr_795  , wr_546  );
  nor g1694( wr_644  , wr_643  , wr_598  );
  nor g1695( wr_559  , wr_558  , wr_530  );
  nor g1696( wr_630  , wr_629  , wr_603  );
  nor g1697( wr_658  , wr_657  , wr_554  );
  nor g1698( wr_974  , wr_973  , wr_863  );
  not g1699( wr_1322 ,           wr_1321 );
  nor g1700( wr_919  , wr_918  , wr_816  );
  nor g1701( wr_1087 , wr_1086 , wr_900  );
  not g1702( wr_2423 ,           wr_2422 );
  not g1703( wr_2444 ,           wr_2443 );
  not g1704( wr_1362 ,           wr_1361 );
  not g1705( wr_1420 ,           wr_1419 );
  nor g1706( wr_2456 , wr_2443 , wr_2422 );
  nor g1707( wr_1010 , wr_1009 , wr_598  );
  nor g1708( wr_1355 , wr_1354 , wr_1351 );
  nor g1709( wr_1364 , wr_1361 , wr_1352 );
  nor g1710( wr_1413 , wr_1412 , wr_1410 );
  nor g1711( wr_1422 , wr_1419 , wr_575  );
  not g1712( wr_2742 ,           wr_2741 );
  not g1713( wr_2772 ,           wr_2771 );
  nor g1714( wr_2797 , wr_2771 , wr_2741 );
  nor g1715( wr_1123 , wr_1122 , wr_530  );
  not g1716( wr_2391 ,           wr_2385 );
  nor g1717( wr_2390 , wr_2389 , wr_2385 );
  not g1718( wr_1041 ,           wr_1040 );
  not g1719( wr_2708 ,           wr_2707 );
  not g1720( wr_2710 ,           wr_2691 );
  not g1721( wr_1154 ,           wr_1153 );
  nor g1722( wr_1277 , wr_1276 , wr_1272 );
  nor g1723( wr_1285 , wr_1284 , wr_1281 );
  not g1724( wr_699  ,           wr_698  );
  not g1725( wr_745  ,           wr_744  );
  nor g1726( wr_702  , wr_698  , wr_701  );
  nor g1727( wr_748  , wr_744  , wr_747  );
  nor g1728( wr_896  , wr_895  , G4091   );
  nor g1729( wr_1002 , wr_1001 , G4091   );
  nor g1730( wr_1058 , wr_1057 , G4091   );
  nor g1731( wr_1835 , wr_1834 , G4091   );
  nor g1732( wr_1848 , wr_1847 , G4091   );
  not g1733( wr_887  ,           wr_886  );
  nor g1734( wr_1180 , wr_1179 , wr_1177 );
  nor g1735( wr_1227 , wr_1226 , wr_1222 );
  nor g1736( wr_1235 , wr_1234 , wr_1231 );
  nor g1737( wr_760  , wr_759  , wr_500  );
  nor g1738( wr_914  , wr_913  , G4091   );
  nor g1739( wr_1115 , wr_1114 , G4091   );
  nor g1740( wr_1147 , wr_1146 , G4091   );
  nor g1741( wr_1171 , wr_1170 , G4091   );
  nor g1742( wr_1191 , wr_1190 , G4091   );
  nor g1743( wr_1877 , wr_1876 , G4091   );
  nor g1744( wr_1890 , wr_1889 , G4091   );
  nor g1745( wr_1903 , wr_1902 , G4091   );
  nor g1746( wr_1916 , wr_1915 , G4091   );
  nor g1747( wr_819  , wr_818  , wr_813  );
  not g1748( wr_905  ,           wr_904  );
  nor g1749( wr_950  , G822    , G4087   );
  nor g1750( wr_1065 , G822    , G4090   );
  nor g1751( wr_1446 , G822    , G1690   );
  nor g1752( wr_1467 , G822    , G1694   );
  not g1753( wr_471  ,           wr_470  );
  nor g1754( wr_513  , wr_512  , wr_484  );
  nor g1755( wr_593  , wr_592  , wr_571  );
  nor g1756( wr_652  , wr_651  , wr_492  );
  not g1757( wr_258  ,           wr_257  );
  not g1758( wr_315  ,           wr_314  );
  not g1759( wr_385  ,           wr_384  );
  nor g1760( wr_938  , wr_937  , wr_576  );
  nor g1761( wr_2217 , wr_2216 , wr_1005 );
  nor g1762( wr_2256 , wr_2255 , wr_979  );
  nor g1763( wr_2269 , wr_2268 , wr_829  );
  nor g1764( wr_2491 , wr_2490 , wr_1118 );
  nor g1765( wr_2543 , wr_2542 , wr_776  );
  not g1766( wr_2208 ,           wr_2207 );
  nor g1767( wr_2307 , wr_2306 , wr_1400 );
  nor g1768( wr_2530 , wr_2529 , wr_1092 );
  nor g1769( wr_1339 , wr_1338 , wr_750  );
  nor g1770( wr_2334 , wr_2333 , wr_816  );
  nor g1771( wr_2481 , wr_1092 , wr_1082 );
  not g1772( wr_2339 ,           wr_2338 );
  nor g1773( wr_2587 , wr_2586 , wr_1314 );
  nor g1774( wr_2614 , wr_2613 , wr_763  );
  not g1775( wr_2619 ,           wr_2618 );
  nor g1776( wr_840  , wr_839  , wr_610  );
  not g1777( wr_788  ,           wr_787  );
  not g1778( wr_645  ,           wr_644  );
  not g1779( wr_560  ,           wr_559  );
  not g1780( wr_631  ,           wr_630  );
  not g1781( wr_659  ,           wr_658  );
  not g1782( wr_975  ,           wr_974  );
  nor g1783( wr_1323 , wr_1322 , wr_763  );
  not g1784( wr_921  ,           wr_919  );
  not g1785( wr_1088 ,           wr_1087 );
  nor g1786( wr_920  , wr_919  , wr_580  );
  nor g1787( wr_2445 , wr_2444 , wr_266  );
  nor g1788( wr_2448 , wr_2443 , wr_2423 );
  nor g1789( wr_2453 , wr_2444 , wr_874  );
  nor g1790( wr_1363 , wr_1362 , wr_508  );
  nor g1791( wr_1421 , wr_1420 , wr_576  );
  not g1792( wr_2457 ,           wr_2456 );
  nor g1793( wr_1014 , wr_1013 , wr_1010 );
  not g1794( wr_1356 ,           wr_1355 );
  not g1795( wr_1414 ,           wr_1413 );
  nor g1796( wr_2785 , wr_2784 , wr_2772 );
  nor g1797( wr_2789 , wr_2771 , wr_2742 );
  nor g1798( wr_2794 , wr_2788 , wr_2772 );
  not g1799( wr_2798 ,           wr_2797 );
  nor g1800( wr_1127 , wr_1126 , wr_1123 );
  nor g1801( wr_2392 , wr_2388 , wr_2391 );
  nor g1802( wr_1042 , wr_1041 , wr_1011 );
  nor g1803( wr_2709 , wr_2708 , wr_2691 );
  nor g1804( wr_2711 , wr_2707 , wr_2710 );
  nor g1805( wr_1155 , wr_1154 , wr_1124 );
  not g1806( wr_1278 ,           wr_1277 );
  not g1807( wr_1286 ,           wr_1285 );
  nor g1808( wr_700  , wr_699  , wr_672  );
  nor g1809( wr_746  , wr_745  , wr_714  );
  nor g1810( wr_897  , wr_896  , wr_892  );
  nor g1811( wr_1003 , wr_1002 , wr_998  );
  nor g1812( wr_1059 , wr_1058 , wr_1054 );
  nor g1813( wr_1836 , wr_1835 , wr_1831 );
  nor g1814( wr_1849 , wr_1848 , wr_1844 );
  nor g1815( wr_888  , wr_887  , wr_861  );
  nor g1816( wr_1181 , wr_1180 , G4092   );
  not g1817( wr_1228 ,           wr_1227 );
  not g1818( wr_1236 ,           wr_1235 );
  nor g1819( wr_766  , wr_765  , wr_760  );
  nor g1820( wr_915  , wr_914  , wr_910  );
  nor g1821( wr_1116 , wr_1115 , wr_1111 );
  nor g1822( wr_1148 , wr_1147 , wr_1143 );
  nor g1823( wr_1172 , wr_1171 , wr_1167 );
  nor g1824( wr_1192 , wr_1191 , wr_1187 );
  nor g1825( wr_1878 , wr_1877 , wr_1873 );
  nor g1826( wr_1891 , wr_1890 , wr_1886 );
  nor g1827( wr_1904 , wr_1903 , wr_1899 );
  nor g1828( wr_1917 , wr_1916 , wr_1912 );
  not g1829( wr_820  ,           wr_819  );
  nor g1830( wr_906  , wr_905  , wr_861  );
  not g1831( wr_951  ,           wr_950  );
  not g1832( wr_1066 ,           wr_1065 );
  not g1833( wr_1447 ,           wr_1446 );
  not g1834( wr_1468 ,           wr_1467 );
  nor g1835( wr_472  , wr_471  , wr_419  );
  not g1836( wr_514  ,           wr_513  );
  not g1837( wr_594  ,           wr_593  );
  not g1838( wr_653  ,           wr_652  );
  nor g1839( wr_259  , wr_258  , wr_217  );
  nor g1840( wr_316  , wr_315  , wr_266  );
  nor g1841( wr_386  , wr_385  , wr_333  );
  not g1842( wr_1293 ,           wr_1180 );
  not g1843( wr_2218 ,           wr_2217 );
  nor g1844( wr_2220 , wr_2217 , wr_597  );
  not g1845( wr_2257 ,           wr_2256 );
  not g1846( wr_2544 ,           wr_2543 );
  not g1847( wr_939  ,           wr_938  );
  not g1848( wr_2270 ,           wr_2269 );
  not g1849( wr_2492 ,           wr_2491 );
  nor g1850( wr_2209 , wr_2208 , wr_825  );
  nor g1851( wr_2308 , wr_2307 , wr_2305 );
  nor g1852( wr_2494 , wr_2491 , wr_782  );
  not g1853( wr_2531 ,           wr_2530 );
  not g1854( wr_1340 ,           wr_1339 );
  not g1855( wr_2335 ,           wr_2334 );
  not g1856( wr_2482 ,           wr_2481 );
  nor g1857( wr_2341 , wr_2338 , wr_2334 );
  nor g1858( wr_2588 , wr_2587 , wr_2585 );
  not g1859( wr_2615 ,           wr_2614 );
  nor g1860( wr_2621 , wr_2618 , wr_2614 );
  nor g1861( wr_848  , wr_847  , wr_840  );
  nor g1862( wr_789  , wr_788  , wr_538  );
  nor g1863( wr_646  , wr_645  , wr_617  );
  nor g1864( wr_561  , wr_560  , wr_522  );
  nor g1865( wr_632  , wr_631  , wr_598  );
  nor g1866( wr_660  , wr_659  , wr_530  );
  nor g1867( wr_976  , wr_975  , wr_598  );
  not g1868( wr_1326 ,           wr_1323 );
  nor g1869( wr_922  , wr_921  , wr_579  );
  nor g1870( wr_1089 , wr_1088 , wr_530  );
  nor g1871( wr_1324 , wr_1323 , wr_500  );
  not g1872( wr_2446 ,           wr_2445 );
  not g1873( wr_2449 ,           wr_2448 );
  not g1874( wr_2454 ,           wr_2453 );
  nor g1875( wr_1365 , wr_1364 , wr_1363 );
  nor g1876( wr_1423 , wr_1422 , wr_1421 );
  nor g1877( wr_2458 , wr_2457 , wr_266  );
  not g1878( wr_1015 ,           wr_1014 );
  not g1879( wr_2786 ,           wr_2785 );
  not g1880( wr_2790 ,           wr_2789 );
  not g1881( wr_2795 ,           wr_2794 );
  nor g1882( wr_2799 , wr_2798 , wr_2784 );
  not g1883( wr_1128 ,           wr_1127 );
  nor g1884( wr_2393 , wr_2392 , wr_2390 );
  not g1885( wr_1043 ,           wr_1042 );
  nor g1886( wr_2712 , wr_2711 , wr_2709 );
  nor g1887( wr_1046 , wr_1042 , wr_1045 );
  not g1888( wr_1156 ,           wr_1155 );
  nor g1889( wr_1287 , wr_1286 , wr_1278 );
  nor g1890( wr_703  , wr_702  , wr_700  );
  nor g1891( wr_749  , wr_748  , wr_746  );
  nor g1892( wr_1159 , wr_1155 , wr_1158 );
  not g1893( wr_898  ,           wr_897  );
  not g1894( wr_1004 ,           wr_1003 );
  not g1895( wr_1060 ,           wr_1059 );
  not g1896( wr_1837 ,           wr_1836 );
  not g1897( wr_1850 ,           wr_1849 );
  not g1898( wr_1182 ,           wr_1181 );
  nor g1899( wr_1237 , wr_1236 , wr_1228 );
  not g1900( wr_767  ,           wr_766  );
  not g1901( wr_916  ,           wr_915  );
  not g1902( wr_1117 ,           wr_1116 );
  not g1903( wr_1149 ,           wr_1148 );
  not g1904( wr_1173 ,           wr_1172 );
  not g1905( wr_1193 ,           wr_1192 );
  not g1906( wr_1879 ,           wr_1878 );
  not g1907( wr_1892 ,           wr_1891 );
  not g1908( wr_1905 ,           wr_1904 );
  not g1909( wr_1918 ,           wr_1917 );
  nor g1910( wr_821  , wr_820  , wr_580  );
  nor g1911( wr_952  , wr_951  , G4088   );
  nor g1912( wr_1067 , wr_1066 , G4089   );
  nor g1913( wr_1448 , wr_1447 , G1689   );
  nor g1914( wr_1469 , wr_1468 , G1691   );
  not g1915( wr_473  ,           wr_472  );
  not g1916( wr_260  ,           wr_259  );
  not g1917( wr_317  ,           wr_316  );
  not g1918( wr_387  ,           wr_386  );
  nor g1919( wr_2219 , wr_2218 , wr_598  );
  nor g1920( wr_2258 , wr_2257 , wr_969  );
  nor g1921( wr_2545 , wr_2544 , wr_1118 );
  nor g1922( wr_940  , wr_939  , wr_816  );
  nor g1923( wr_2271 , wr_2270 , wr_1005 );
  nor g1924( wr_2493 , wr_2492 , wr_781  );
  not g1925( wr_2210 ,           wr_2209 );
  not g1926( wr_2309 ,           wr_2308 );
  nor g1927( wr_2532 , wr_2531 , wr_1082 );
  nor g1928( wr_1341 , wr_1340 , wr_763  );
  nor g1929( wr_2340 , wr_2339 , wr_2335 );
  nor g1930( wr_2483 , wr_2482 , wr_772  );
  not g1931( wr_2589 ,           wr_2588 );
  nor g1932( wr_2620 , wr_2619 , wr_2615 );
  not g1933( wr_849  ,           wr_848  );
  nor g1934( wr_797  , wr_796  , wr_789  );
  not g1935( wr_633  ,           wr_632  );
  not g1936( wr_661  ,           wr_660  );
  nor g1937( wr_980  , wr_979  , wr_976  );
  nor g1938( wr_1327 , wr_1326 , wr_1325 );
  nor g1939( wr_923  , wr_922  , wr_920  );
  nor g1940( wr_1093 , wr_1092 , wr_1089 );
  nor g1941( wr_2447 , wr_2446 , wr_2423 );
  nor g1942( wr_2450 , wr_2449 , wr_874  );
  nor g1943( wr_2455 , wr_2454 , wr_2422 );
  nor g1944( wr_1016 , wr_1015 , wr_829  );
  nor g1945( wr_2787 , wr_2786 , wr_2742 );
  nor g1946( wr_2791 , wr_2790 , wr_2788 );
  nor g1947( wr_2796 , wr_2795 , wr_2741 );
  nor g1948( wr_1129 , wr_1128 , wr_776  );
  not g1949( wr_2464 ,           wr_2393 );
  nor g1950( wr_1044 , wr_1043 , wr_610  );
  not g1951( wr_2805 ,           wr_2712 );
  nor g1952( wr_1157 , wr_1156 , wr_538  );
  not g1953( wr_1288 ,           wr_1287 );
  not g1954( G1002   ,           wr_703  );
  not g1955( G1004   ,           wr_749  );
  nor g1956( wr_1291 , wr_1287 , wr_1290 );
  nor g1957( G838    , wr_898  , wr_888  );
  nor g1958( wr_1183 , wr_1182 , wr_861  );
  not g1959( wr_1238 ,           wr_1237 );
  nor g1960( wr_768  , wr_767  , wr_753  );
  nor g1961( G861    , wr_916  , wr_906  );
  nor g1962( wr_1241 , wr_1237 , wr_1240 );
  not g1963( wr_822  ,           wr_821  );
  nor g1964( wr_964  , wr_963  , wr_952  );
  nor g1965( wr_1077 , wr_1076 , wr_1067 );
  nor g1966( wr_1460 , wr_1459 , wr_1448 );
  nor g1967( wr_1479 , wr_1478 , wr_1469 );
  nor g1968( wr_474  , wr_473  , wr_403  );
  not g1969( wr_562  ,           wr_561  );
  not g1970( wr_647  ,           wr_646  );
  nor g1971( G598    , wr_317  , wr_260  );
  nor g1972( wr_2221 , wr_2220 , wr_2219 );
  not g1973( wr_2259 ,           wr_2258 );
  not g1974( wr_2548 ,           wr_2545 );
  not g1975( wr_941  ,           wr_940  );
  not g1976( wr_2272 ,           wr_2271 );
  nor g1977( wr_2495 , wr_2494 , wr_2493 );
  nor g1978( wr_2547 , wr_2546 , wr_2545 );
  nor g1979( wr_2211 , wr_2210 , wr_831  );
  nor g1980( wr_2275 , wr_2271 , wr_2274 );
  nor g1981( wr_2310 , wr_2309 , wr_940  );
  not g1982( wr_2533 ,           wr_2532 );
  not g1983( wr_1342 ,           wr_1341 );
  nor g1984( wr_2342 , wr_2341 , wr_2340 );
  not g1985( wr_2484 ,           wr_2483 );
  nor g1986( wr_2590 , wr_2589 , wr_1341 );
  nor g1987( wr_2622 , wr_2621 , wr_2620 );
  nor g1988( wr_850  , wr_849  , wr_833  );
  not g1989( wr_798  ,           wr_797  );
  nor g1990( wr_926  , wr_633  , wr_863  );
  nor g1991( wr_1299 , wr_661  , wr_900  );
  nor g1992( wr_943  , wr_940  , wr_579  );
  not g1993( wr_981  ,           wr_980  );
  nor g1994( wr_1328 , wr_1327 , wr_1324 );
  nor g1995( wr_1344 , wr_1341 , wr_1325 );
  not g1996( wr_924  ,           wr_923  );
  not g1997( wr_1094 ,           wr_1093 );
  nor g1998( wr_2451 , wr_2450 , wr_2447 );
  nor g1999( wr_2459 , wr_2458 , wr_2455 );
  not g2000( wr_1017 ,           wr_1016 );
  nor g2001( wr_2792 , wr_2791 , wr_2787 );
  nor g2002( wr_2800 , wr_2799 , wr_2796 );
  not g2003( wr_1130 ,           wr_1129 );
  nor g2004( wr_1047 , wr_1046 , wr_1044 );
  nor g2005( wr_1160 , wr_1159 , wr_1157 );
  nor g2006( wr_1289 , wr_1288 , wr_1253 );
  nor g2007( wr_1851 , G1004   , G1002   );
  nor g2008( wr_1542 , G838    , G4087   );
  nor g2009( wr_1612 , G838    , G4090   );
  nor g2010( wr_1648 , G838    , G1690   );
  nor g2011( wr_1722 , G838    , G1694   );
  nor g2012( G877    , wr_1193 , wr_1183 );
  nor g2013( wr_1239 , wr_1238 , wr_1203 );
  not g2014( wr_769  ,           wr_768  );
  nor g2015( wr_947  , G861    , G4087   );
  nor g2016( wr_1062 , G861    , G4090   );
  nor g2017( wr_1443 , G861    , G1690   );
  nor g2018( wr_1464 , G861    , G1694   );
  nor g2019( wr_823  , wr_822  , wr_806  );
  not g2020( wr_965  ,           wr_964  );
  not g2021( wr_1078 ,           wr_1077 );
  not g2022( wr_1461 ,           wr_1460 );
  not g2023( wr_1480 ,           wr_1479 );
  not g2024( wr_475  ,           wr_474  );
  nor g2025( G588    , wr_562  , wr_514  );
  nor g2026( G615    , wr_633  , wr_594  );
  nor g2027( G626    , wr_647  , wr_639  );
  nor g2028( G632    , wr_661  , wr_653  );
  not g2029( wr_2222 ,           wr_2221 );
  nor g2030( wr_2224 , wr_2221 , wr_2213 );
  nor g2031( wr_2260 , wr_2259 , wr_825  );
  nor g2032( wr_2550 , wr_2549 , wr_2548 );
  nor g2033( wr_2273 , wr_2272 , wr_2264 );
  nor g2034( wr_2311 , wr_2308 , wr_941  );
  not g2035( wr_2496 ,           wr_2495 );
  not g2036( wr_2212 ,           wr_2211 );
  nor g2037( wr_2498 , wr_2495 , wr_2487 );
  nor g2038( wr_2534 , wr_2533 , wr_772  );
  not g2039( wr_2343 ,           wr_2342 );
  nor g2040( wr_2485 , wr_2484 , wr_778  );
  nor g2041( wr_2591 , wr_2588 , wr_1342 );
  nor g2042( wr_2345 , wr_2342 , wr_1389 );
  not g2043( wr_2623 ,           wr_2622 );
  nor g2044( wr_2625 , wr_2622 , wr_1303 );
  not g2045( wr_851  ,           wr_850  );
  nor g2046( wr_799  , wr_798  , wr_780  );
  nor g2047( wr_942  , wr_941  , wr_580  );
  nor g2048( wr_1343 , wr_1342 , wr_500  );
  nor g2049( wr_982  , wr_981  , wr_969  );
  not g2050( wr_1329 ,           wr_1328 );
  nor g2051( wr_1095 , wr_1094 , wr_1082 );
  not g2052( wr_2452 ,           wr_2451 );
  not g2053( wr_2460 ,           wr_2459 );
  nor g2054( wr_1018 , wr_1017 , wr_1005 );
  not g2055( wr_2793 ,           wr_2792 );
  not g2056( wr_2801 ,           wr_2800 );
  nor g2057( wr_1131 , wr_1130 , wr_1118 );
  nor g2058( wr_1048 , wr_1047 , G4092   );
  nor g2059( wr_1161 , wr_1160 , G4092   );
  nor g2060( wr_1292 , wr_1291 , wr_1289 );
  not g2061( wr_1852 ,           wr_1851 );
  not g2062( wr_1295 ,           wr_1160 );
  not g2063( wr_1385 ,           wr_1047 );
  not g2064( wr_1543 ,           wr_1542 );
  not g2065( wr_1613 ,           wr_1612 );
  not g2066( wr_1649 ,           wr_1648 );
  not g2067( wr_1723 ,           wr_1722 );
  nor g2068( wr_1242 , wr_1241 , wr_1239 );
  nor g2069( wr_1539 , G877    , G4087   );
  nor g2070( wr_1609 , G877    , G4090   );
  nor g2071( wr_1645 , G877    , G1690   );
  nor g2072( wr_1719 , G877    , G1694   );
  nor g2073( wr_770  , wr_769  , wr_752  );
  not g2074( wr_948  ,           wr_947  );
  not g2075( wr_1063 ,           wr_1062 );
  not g2076( wr_1444 ,           wr_1443 );
  not g2077( wr_1465 ,           wr_1464 );
  not g2078( wr_824  ,           wr_823  );
  nor g2079( G610    , wr_475  , wr_387  );
  nor g2080( wr_2223 , wr_2222 , wr_2214 );
  not g2081( wr_2261 ,           wr_2260 );
  nor g2082( wr_2551 , wr_2550 , wr_2547 );
  nor g2083( wr_2276 , wr_2275 , wr_2273 );
  nor g2084( wr_2312 , wr_2311 , wr_2310 );
  nor g2085( wr_2497 , wr_2496 , wr_2488 );
  not g2086( wr_2535 ,           wr_2534 );
  nor g2087( wr_2344 , wr_2343 , wr_571  );
  not g2088( wr_2486 ,           wr_2485 );
  nor g2089( wr_2592 , wr_2591 , wr_2590 );
  nor g2090( wr_2624 , wr_2623 , wr_492  );
  nor g2091( wr_852  , wr_851  , wr_828  );
  not g2092( wr_800  ,           wr_799  );
  nor g2093( wr_944  , wr_943  , wr_942  );
  nor g2094( wr_1345 , wr_1344 , wr_1343 );
  not g2095( wr_983  ,           wr_982  );
  not g2096( wr_1096 ,           wr_1095 );
  nor g2097( wr_2461 , wr_2460 , wr_2452 );
  not g2098( wr_1019 ,           wr_1018 );
  nor g2099( wr_2802 , wr_2801 , wr_2793 );
  nor g2100( wr_1022 , wr_1018 , wr_1021 );
  not g2101( wr_1132 ,           wr_1131 );
  nor g2102( wr_1135 , wr_1131 , wr_1134 );
  not g2103( wr_1049 ,           wr_1048 );
  not g2104( wr_1162 ,           wr_1161 );
  not g2105( G1000   ,           wr_1292 );
  nor g2106( wr_1544 , wr_1543 , G4088   );
  nor g2107( wr_1614 , wr_1613 , G4089   );
  nor g2108( wr_1650 , wr_1649 , G1689   );
  nor g2109( wr_1724 , wr_1723 , G1691   );
  not g2110( G998    ,           wr_1242 );
  not g2111( wr_1540 ,           wr_1539 );
  not g2112( wr_1610 ,           wr_1609 );
  not g2113( wr_1646 ,           wr_1645 );
  not g2114( wr_1720 ,           wr_1719 );
  not g2115( wr_771  ,           wr_770  );
  nor g2116( wr_949  , wr_948  , wr_946  );
  nor g2117( wr_1064 , wr_1063 , wr_1061 );
  nor g2118( wr_1445 , wr_1444 , wr_1442 );
  nor g2119( wr_1466 , wr_1465 , wr_1463 );
  nor g2120( wr_2225 , wr_2224 , wr_2223 );
  nor g2121( wr_2262 , wr_2261 , wr_831  );
  not g2122( wr_2552 ,           wr_2551 );
  not g2123( wr_2277 ,           wr_2276 );
  not g2124( wr_2313 ,           wr_2312 );
  nor g2125( wr_2499 , wr_2498 , wr_2497 );
  nor g2126( wr_2555 , wr_2551 , wr_2554 );
  nor g2127( wr_2315 , wr_2312 , wr_1389 );
  nor g2128( wr_2536 , wr_2535 , wr_778  );
  nor g2129( wr_2346 , wr_2345 , wr_2344 );
  not g2130( wr_2593 ,           wr_2592 );
  nor g2131( wr_2595 , wr_2592 , wr_1303 );
  nor g2132( wr_2626 , wr_2625 , wr_2624 );
  not g2133( wr_853  ,           wr_852  );
  nor g2134( wr_801  , wr_800  , wr_775  );
  nor g2135( wr_984  , wr_983  , wr_825  );
  nor g2136( wr_1097 , wr_1096 , wr_772  );
  not g2137( wr_2462 ,           wr_2461 );
  nor g2138( wr_2465 , wr_2461 , wr_2464 );
  nor g2139( wr_1020 , wr_1019 , wr_603  );
  not g2140( wr_2803 ,           wr_2802 );
  nor g2141( wr_2806 , wr_2802 , wr_2805 );
  nor g2142( wr_1133 , wr_1132 , wr_554  );
  nor g2143( wr_1050 , wr_1049 , wr_861  );
  nor g2144( wr_1163 , wr_1162 , wr_861  );
  nor g2145( wr_1853 , wr_1852 , G1000   );
  nor g2146( wr_1555 , wr_1554 , wr_1544 );
  nor g2147( wr_1623 , wr_1622 , wr_1614 );
  nor g2148( wr_1661 , wr_1660 , wr_1650 );
  nor g2149( wr_1733 , wr_1732 , wr_1724 );
  nor g2150( wr_1541 , wr_1540 , wr_946  );
  nor g2151( wr_1611 , wr_1610 , wr_1061 );
  nor g2152( wr_1647 , wr_1646 , wr_1442 );
  nor g2153( wr_1721 , wr_1720 , wr_1463 );
  nor g2154( wr_966  , wr_965  , wr_949  );
  nor g2155( wr_1079 , wr_1078 , wr_1064 );
  nor g2156( wr_1462 , wr_1461 , wr_1445 );
  nor g2157( wr_1481 , wr_1480 , wr_1466 );
  not g2158( wr_2226 ,           wr_2225 );
  nor g2159( wr_2228 , wr_2225 , wr_2211 );
  not g2160( wr_2279 ,           wr_2262 );
  nor g2161( wr_2553 , wr_2552 , wr_2538 );
  nor g2162( wr_2278 , wr_2277 , wr_2262 );
  nor g2163( wr_2314 , wr_2313 , wr_571  );
  not g2164( wr_2500 ,           wr_2499 );
  nor g2165( wr_2502 , wr_2499 , wr_2485 );
  not g2166( wr_2559 ,           wr_2536 );
  not g2167( wr_2347 ,           wr_2346 );
  nor g2168( wr_2594 , wr_2593 , wr_492  );
  nor g2169( wr_2349 , wr_2346 , wr_1394 );
  not g2170( wr_2627 ,           wr_2626 );
  nor g2171( wr_2629 , wr_2626 , wr_1308 );
  nor g2172( wr_854  , wr_853  , wr_827  );
  not g2173( wr_802  ,           wr_801  );
  not g2174( wr_985  ,           wr_984  );
  not g2175( wr_1098 ,           wr_1097 );
  nor g2176( wr_2463 , wr_2462 , wr_2393 );
  nor g2177( wr_1023 , wr_1022 , wr_1020 );
  nor g2178( wr_2804 , wr_2803 , wr_2712 );
  nor g2179( wr_1136 , wr_1135 , wr_1133 );
  nor g2180( G836    , wr_1060 , wr_1050 );
  nor g2181( G875    , wr_1173 , wr_1163 );
  not g2182( wr_1854 ,           wr_1853 );
  not g2183( wr_1556 ,           wr_1555 );
  not g2184( wr_1624 ,           wr_1623 );
  not g2185( wr_1662 ,           wr_1661 );
  not g2186( wr_1734 ,           wr_1733 );
  not g2187( G722    ,           wr_966  );
  not g2188( G859    ,           wr_1079 );
  nor g2189( G661    , wr_1462 , wr_1441 );
  nor g2190( G693    , wr_1481 , wr_1441 );
  nor g2191( wr_2227 , wr_2226 , wr_2212 );
  nor g2192( wr_2280 , wr_2276 , wr_2279 );
  nor g2193( wr_2556 , wr_2555 , wr_2553 );
  nor g2194( wr_2316 , wr_2315 , wr_2314 );
  nor g2195( wr_2501 , wr_2500 , wr_2486 );
  nor g2196( wr_2348 , wr_2347 , wr_588  );
  nor g2197( wr_2596 , wr_2595 , wr_2594 );
  nor g2198( wr_2628 , wr_2627 , wr_484  );
  not g2199( wr_925  ,           wr_854  );
  nor g2200( wr_803  , wr_802  , wr_774  );
  nor g2201( wr_986  , wr_985  , wr_831  );
  nor g2202( wr_1099 , wr_1098 , wr_778  );
  nor g2203( wr_2466 , wr_2465 , wr_2463 );
  nor g2204( wr_1024 , wr_1023 , G4092   );
  nor g2205( wr_2807 , wr_2806 , wr_2804 );
  nor g2206( wr_1137 , wr_1136 , G4092   );
  not g2207( wr_1296 ,           wr_1136 );
  not g2208( wr_1386 ,           wr_1023 );
  nor g2209( wr_1523 , G836    , G4087   );
  nor g2210( wr_1595 , G836    , G4090   );
  nor g2211( wr_1667 , G836    , G1690   );
  nor g2212( wr_1739 , G836    , G1694   );
  nor g2213( wr_1520 , G875    , G4087   );
  nor g2214( wr_1592 , G875    , G4090   );
  nor g2215( wr_1664 , G875    , G1690   );
  nor g2216( wr_1736 , G875    , G1694   );
  nor g2217( wr_1855 , wr_1854 , G850    );
  nor g2218( wr_855  , wr_854  , wr_594  );
  nor g2219( wr_859  , wr_854  , wr_639  );
  nor g2220( wr_1557 , wr_1556 , wr_1541 );
  nor g2221( wr_1625 , wr_1624 , wr_1611 );
  nor g2222( wr_1663 , wr_1662 , wr_1647 );
  nor g2223( wr_1735 , wr_1734 , wr_1721 );
  nor g2224( wr_2229 , wr_2228 , wr_2227 );
  nor g2225( wr_2281 , wr_2280 , wr_2278 );
  not g2226( wr_2557 ,           wr_2556 );
  not g2227( wr_2317 ,           wr_2316 );
  nor g2228( wr_2503 , wr_2502 , wr_2501 );
  nor g2229( wr_2560 , wr_2556 , wr_2559 );
  nor g2230( wr_2319 , wr_2316 , wr_1394 );
  nor g2231( wr_2350 , wr_2349 , wr_2348 );
  not g2232( wr_2597 ,           wr_2596 );
  nor g2233( wr_2599 , wr_2596 , wr_1308 );
  nor g2234( wr_2630 , wr_2629 , wr_2628 );
  nor g2235( wr_2362 , wr_925  , wr_646  );
  not g2236( wr_1298 ,           wr_803  );
  nor g2237( wr_927  , wr_926  , wr_925  );
  not g2238( wr_987  ,           wr_986  );
  nor g2239( wr_990  , wr_986  , wr_989  );
  not g2240( wr_1100 ,           wr_1099 );
  nor g2241( wr_1103 , wr_1099 , wr_1102 );
  nor g2242( wr_2832 , wr_2466 , G4091   );
  not g2243( wr_1025 ,           wr_1024 );
  nor g2244( wr_2821 , wr_2807 , G4091   );
  not g2245( wr_1138 ,           wr_1137 );
  not g2246( wr_2467 ,           wr_2466 );
  not g2247( wr_2808 ,           wr_2807 );
  not g2248( wr_1524 ,           wr_1523 );
  not g2249( wr_1596 ,           wr_1595 );
  not g2250( wr_1668 ,           wr_1667 );
  not g2251( wr_1740 ,           wr_1739 );
  not g2252( wr_1521 ,           wr_1520 );
  not g2253( wr_1593 ,           wr_1592 );
  not g2254( wr_1665 ,           wr_1664 );
  not g2255( wr_1737 ,           wr_1736 );
  not g2256( wr_1856 ,           wr_1855 );
  nor g2257( wr_804  , wr_803  , wr_514  );
  nor g2258( wr_857  , wr_803  , wr_653  );
  nor g2259( wr_856  , wr_855  , wr_824  );
  nor g2260( wr_860  , wr_859  , wr_824  );
  not g2261( G762    ,           wr_1557 );
  not g2262( G802    ,           wr_1625 );
  nor g2263( G664    , wr_1663 , wr_1441 );
  nor g2264( G696    , wr_1735 , wr_1441 );
  not g2265( wr_2230 ,           wr_2229 );
  nor g2266( wr_2232 , wr_2229 , wr_597  );
  not g2267( wr_2282 ,           wr_2281 );
  nor g2268( wr_2558 , wr_2557 , wr_2536 );
  nor g2269( wr_2284 , wr_2281 , wr_597  );
  nor g2270( wr_2318 , wr_2317 , wr_588  );
  not g2271( wr_2504 ,           wr_2503 );
  nor g2272( wr_2506 , wr_2503 , wr_901  );
  not g2273( wr_2351 ,           wr_2350 );
  nor g2274( wr_2598 , wr_2597 , wr_484  );
  nor g2275( wr_2353 , wr_2350 , wr_579  );
  not g2276( wr_2631 ,           wr_2630 );
  nor g2277( wr_2633 , wr_2630 , wr_1325 );
  not g2278( wr_2366 ,           wr_2362 );
  nor g2279( wr_2642 , wr_1298 , wr_561  );
  nor g2280( wr_1300 , wr_1299 , wr_1298 );
  not g2281( wr_928  ,           wr_927  );
  nor g2282( wr_945  , wr_944  , wr_927  );
  nor g2283( wr_1424 , wr_1423 , wr_927  );
  nor g2284( wr_1404 , wr_1403 , wr_927  );
  nor g2285( wr_1390 , wr_927  , wr_1389 );
  nor g2286( wr_988  , wr_987  , wr_625  );
  nor g2287( wr_1101 , wr_1100 , wr_546  );
  nor g2288( wr_1026 , wr_1025 , wr_861  );
  nor g2289( wr_1139 , wr_1138 , wr_861  );
  nor g2290( wr_2468 , wr_2467 , G4092   );
  nor g2291( wr_2809 , wr_2808 , G4092   );
  nor g2292( wr_1525 , wr_1524 , G4088   );
  nor g2293( wr_1597 , wr_1596 , G4089   );
  nor g2294( wr_1669 , wr_1668 , G1689   );
  nor g2295( wr_1741 , wr_1740 , G1691   );
  nor g2296( wr_1522 , wr_1521 , wr_946  );
  nor g2297( wr_1594 , wr_1593 , wr_1061 );
  nor g2298( wr_1666 , wr_1665 , wr_1442 );
  nor g2299( wr_1738 , wr_1737 , wr_1463 );
  nor g2300( wr_1857 , wr_1856 , G998    );
  nor g2301( wr_805  , wr_804  , wr_771  );
  nor g2302( wr_858  , wr_857  , wr_771  );
  not g2303( G618    ,           wr_856  );
  not g2304( G629    ,           wr_860  );
  nor g2305( wr_2231 , wr_2230 , wr_598  );
  nor g2306( wr_2283 , wr_2282 , wr_598  );
  nor g2307( wr_2561 , wr_2560 , wr_2558 );
  nor g2308( wr_2320 , wr_2319 , wr_2318 );
  nor g2309( wr_2505 , wr_2504 , wr_530  );
  nor g2310( wr_2352 , wr_2351 , wr_580  );
  nor g2311( wr_2600 , wr_2599 , wr_2598 );
  nor g2312( wr_2632 , wr_2631 , wr_500  );
  not g2313( wr_2646 ,           wr_2642 );
  not g2314( wr_1301 ,           wr_1300 );
  nor g2315( wr_929  , wr_928  , wr_924  );
  nor g2316( wr_1346 , wr_1345 , wr_1300 );
  nor g2317( wr_1366 , wr_1365 , wr_1300 );
  nor g2318( wr_1415 , wr_1414 , wr_928  );
  nor g2319( wr_1318 , wr_1317 , wr_1300 );
  nor g2320( wr_1397 , wr_1396 , wr_928  );
  nor g2321( wr_1304 , wr_1300 , wr_1303 );
  nor g2322( wr_1388 , wr_928  , wr_571  );
  nor g2323( wr_991  , wr_990  , wr_988  );
  nor g2324( wr_1104 , wr_1103 , wr_1101 );
  nor g2325( G834    , wr_1036 , wr_1026 );
  nor g2326( G873    , wr_1149 , wr_1139 );
  not g2327( wr_2469 ,           wr_2468 );
  not g2328( wr_2810 ,           wr_2809 );
  nor g2329( wr_1536 , wr_1535 , wr_1525 );
  nor g2330( wr_1606 , wr_1605 , wr_1597 );
  nor g2331( wr_1680 , wr_1679 , wr_1669 );
  nor g2332( wr_1750 , wr_1749 , wr_1741 );
  not g2333( wr_1858 ,           wr_1857 );
  not g2334( G591    ,           wr_805  );
  not g2335( G621    ,           wr_858  );
  nor g2336( wr_2233 , wr_2232 , wr_2231 );
  nor g2337( wr_2285 , wr_2284 , wr_2283 );
  not g2338( wr_2562 ,           wr_2561 );
  not g2339( wr_2321 ,           wr_2320 );
  nor g2340( wr_2507 , wr_2506 , wr_2505 );
  nor g2341( wr_2564 , wr_2561 , wr_901  );
  nor g2342( wr_2323 , wr_2320 , wr_579  );
  nor g2343( wr_2354 , wr_2353 , wr_2352 );
  not g2344( wr_2601 ,           wr_2600 );
  nor g2345( wr_2603 , wr_2600 , wr_1325 );
  nor g2346( wr_2634 , wr_2633 , wr_2632 );
  nor g2347( wr_1330 , wr_1329 , wr_1301 );
  nor g2348( wr_1357 , wr_1356 , wr_1301 );
  nor g2349( G623    , wr_945  , wr_929  );
  nor g2350( wr_1425 , wr_1424 , wr_1415 );
  nor g2351( wr_1311 , wr_1310 , wr_1301 );
  nor g2352( wr_1405 , wr_1404 , wr_1397 );
  nor g2353( wr_1302 , wr_1301 , wr_492  );
  nor g2354( wr_1391 , wr_1390 , wr_1388 );
  nor g2355( wr_992  , wr_991  , G4092   );
  not g2356( wr_1297 ,           wr_1104 );
  not g2357( wr_1387 ,           wr_991  );
  nor g2358( wr_1105 , wr_1104 , G4092   );
  nor g2359( wr_1504 , G834    , G4087   );
  nor g2360( wr_1578 , G834    , G4090   );
  nor g2361( wr_1686 , G834    , G1690   );
  nor g2362( wr_1756 , G834    , G1694   );
  nor g2363( wr_1501 , G873    , G4087   );
  nor g2364( wr_1575 , G873    , G4090   );
  nor g2365( wr_1683 , G873    , G1690   );
  nor g2366( wr_1753 , G873    , G1694   );
  nor g2367( wr_2470 , wr_2469 , G4091   );
  nor g2368( wr_2811 , wr_2810 , G4091   );
  not g2369( wr_1537 ,           wr_1536 );
  not g2370( wr_1607 ,           wr_1606 );
  not g2371( wr_1681 ,           wr_1680 );
  not g2372( wr_1751 ,           wr_1750 );
  nor g2373( G854    , wr_1866 , wr_1858 );
  not g2374( wr_2234 ,           wr_2233 );
  nor g2375( wr_2236 , wr_2233 , wr_883  );
  not g2376( wr_2286 ,           wr_2285 );
  nor g2377( wr_2563 , wr_2562 , wr_530  );
  nor g2378( wr_2288 , wr_2285 , wr_883  );
  nor g2379( wr_2322 , wr_2321 , wr_580  );
  not g2380( wr_2508 ,           wr_2507 );
  nor g2381( wr_2510 , wr_2507 , wr_1178 );
  not g2382( wr_2355 ,           wr_2354 );
  nor g2383( wr_2602 , wr_2601 , wr_500  );
  nor g2384( wr_2357 , wr_2354 , wr_575  );
  not g2385( wr_2635 ,           wr_2634 );
  nor g2386( wr_2637 , wr_2634 , wr_1352 );
  nor g2387( wr_1347 , wr_1346 , wr_1330 );
  nor g2388( wr_1367 , wr_1366 , wr_1357 );
  not g2389( wr_1407 ,           G623    );
  not g2390( wr_1426 ,           wr_1425 );
  nor g2391( wr_1319 , wr_1318 , wr_1311 );
  not g2392( wr_1406 ,           wr_1405 );
  nor g2393( wr_1305 , wr_1304 , wr_1302 );
  not g2394( wr_1392 ,           wr_1391 );
  nor g2395( wr_1801 , G623    , G4092   );
  nor g2396( wr_1812 , wr_1425 , G4092   );
  nor g2397( wr_1825 , wr_1405 , G4092   );
  nor g2398( wr_1838 , wr_1391 , G4092   );
  not g2399( wr_993  ,           wr_992  );
  nor g2400( wr_1785 , G623    , wr_1784 );
  not g2401( wr_1106 ,           wr_1105 );
  not g2402( wr_1505 ,           wr_1504 );
  not g2403( wr_1579 ,           wr_1578 );
  not g2404( wr_1687 ,           wr_1686 );
  not g2405( wr_1757 ,           wr_1756 );
  not g2406( wr_1502 ,           wr_1501 );
  not g2407( wr_1576 ,           wr_1575 );
  not g2408( wr_1684 ,           wr_1683 );
  not g2409( wr_1754 ,           wr_1753 );
  nor g2410( wr_2478 , wr_2477 , wr_2470 );
  nor g2411( wr_2818 , wr_2817 , wr_2811 );
  nor g2412( wr_1799 , wr_1798 , G623    );
  nor g2413( wr_1538 , wr_1537 , wr_1522 );
  nor g2414( wr_1608 , wr_1607 , wr_1594 );
  nor g2415( wr_1682 , wr_1681 , wr_1666 );
  nor g2416( wr_1752 , wr_1751 , wr_1738 );
  nor g2417( wr_2235 , wr_2234 , wr_617  );
  nor g2418( wr_2287 , wr_2286 , wr_617  );
  nor g2419( wr_2565 , wr_2564 , wr_2563 );
  nor g2420( wr_2324 , wr_2323 , wr_2322 );
  nor g2421( wr_2509 , wr_2508 , wr_522  );
  nor g2422( wr_2356 , wr_2355 , wr_576  );
  nor g2423( wr_2604 , wr_2603 , wr_2602 );
  nor g2424( wr_2636 , wr_2635 , wr_508  );
  not g2425( wr_1348 ,           wr_1347 );
  not g2426( wr_1368 ,           wr_1367 );
  nor g2427( wr_1427 , wr_1426 , wr_1407 );
  not g2428( wr_1320 ,           wr_1319 );
  not g2429( wr_1306 ,           wr_1305 );
  not g2430( wr_1802 ,           wr_1801 );
  not g2431( wr_1813 ,           wr_1812 );
  not g2432( wr_1826 ,           wr_1825 );
  not g2433( wr_1839 ,           wr_1838 );
  nor g2434( wr_994  , wr_993  , wr_861  );
  nor g2435( wr_1867 , wr_1347 , G4092   );
  nor g2436( wr_1880 , wr_1367 , G4092   );
  nor g2437( wr_1893 , wr_1319 , G4092   );
  nor g2438( wr_1906 , wr_1305 , G4092   );
  not g2439( wr_1786 ,           wr_1785 );
  nor g2440( wr_1107 , wr_1106 , wr_861  );
  nor g2441( wr_1506 , wr_1505 , G4088   );
  nor g2442( wr_1580 , wr_1579 , G4089   );
  nor g2443( wr_1688 , wr_1687 , G1689   );
  nor g2444( wr_1758 , wr_1757 , G1691   );
  nor g2445( wr_1503 , wr_1502 , wr_946  );
  nor g2446( wr_1577 , wr_1576 , wr_1061 );
  nor g2447( wr_1685 , wr_1684 , wr_1442 );
  nor g2448( wr_1755 , wr_1754 , wr_1463 );
  nor g2449( wr_1797 , wr_1777 , wr_1407 );
  not g2450( wr_2479 ,           wr_2478 );
  not g2451( wr_2819 ,           wr_2818 );
  not g2452( G757    ,           wr_1538 );
  not g2453( G797    ,           wr_1608 );
  nor g2454( G667    , wr_1682 , wr_1441 );
  nor g2455( G699    , wr_1752 , wr_1441 );
  nor g2456( wr_2237 , wr_2236 , wr_2235 );
  nor g2457( wr_2289 , wr_2288 , wr_2287 );
  not g2458( wr_2566 ,           wr_2565 );
  not g2459( wr_2325 ,           wr_2324 );
  nor g2460( wr_2511 , wr_2510 , wr_2509 );
  nor g2461( wr_2568 , wr_2565 , wr_1178 );
  nor g2462( wr_2327 , wr_2324 , wr_575  );
  nor g2463( wr_2358 , wr_2357 , wr_2356 );
  not g2464( wr_2605 ,           wr_2604 );
  nor g2465( wr_2607 , wr_2604 , wr_1352 );
  nor g2466( wr_2638 , wr_2637 , wr_2636 );
  nor g2467( wr_1369 , wr_1368 , wr_1348 );
  not g2468( wr_1428 ,           wr_1427 );
  nor g2469( wr_1803 , wr_1802 , wr_861  );
  nor g2470( wr_1814 , wr_1813 , wr_861  );
  nor g2471( wr_1827 , wr_1826 , wr_861  );
  nor g2472( wr_1840 , wr_1839 , wr_861  );
  nor g2473( G832    , wr_1004 , wr_994  );
  not g2474( wr_1868 ,           wr_1867 );
  not g2475( wr_1881 ,           wr_1880 );
  not g2476( wr_1894 ,           wr_1893 );
  not g2477( wr_1907 ,           wr_1906 );
  nor g2478( wr_1787 , wr_1786 , wr_1773 );
  nor g2479( G871    , wr_1117 , wr_1107 );
  nor g2480( wr_1517 , wr_1516 , wr_1506 );
  nor g2481( wr_1589 , wr_1588 , wr_1580 );
  nor g2482( wr_1699 , wr_1698 , wr_1688 );
  nor g2483( wr_1767 , wr_1766 , wr_1758 );
  nor g2484( wr_1800 , wr_1799 , wr_1797 );
  not g2485( wr_2238 ,           wr_2237 );
  nor g2486( wr_2240 , wr_2237 , wr_989  );
  not g2487( wr_2290 ,           wr_2289 );
  nor g2488( wr_2567 , wr_2566 , wr_522  );
  nor g2489( wr_2292 , wr_2289 , wr_989  );
  nor g2490( wr_2326 , wr_2325 , wr_576  );
  not g2491( wr_2512 ,           wr_2511 );
  nor g2492( wr_2514 , wr_2511 , wr_1102 );
  nor g2493( wr_2367 , wr_2358 , wr_2252 );
  nor g2494( wr_2606 , wr_2605 , wr_508  );
  nor g2495( wr_2359 , wr_2358 , G2174   );
  nor g2496( wr_2647 , wr_2638 , wr_2526 );
  nor g2497( wr_2639 , wr_2638 , G1497   );
  not g2498( wr_1370 ,           wr_1369 );
  nor g2499( wr_1429 , wr_1428 , wr_1406 );
  nor g2500( G824    , wr_1811 , wr_1803 );
  nor g2501( G826    , wr_1824 , wr_1814 );
  nor g2502( G828    , wr_1837 , wr_1827 );
  nor g2503( G830    , wr_1850 , wr_1840 );
  nor g2504( wr_1485 , G832    , G4087   );
  nor g2505( wr_1561 , G832    , G4090   );
  nor g2506( wr_1629 , G832    , G1690   );
  nor g2507( wr_1705 , G832    , G1694   );
  nor g2508( wr_1869 , wr_1868 , wr_861  );
  nor g2509( wr_1882 , wr_1881 , wr_861  );
  nor g2510( wr_1895 , wr_1894 , wr_861  );
  nor g2511( wr_1908 , wr_1907 , wr_861  );
  nor g2512( wr_1792 , wr_1791 , wr_1787 );
  nor g2513( wr_1482 , G871    , G4087   );
  nor g2514( wr_1558 , G871    , G4090   );
  nor g2515( wr_1626 , G871    , G1690   );
  nor g2516( wr_1702 , G871    , G1694   );
  not g2517( wr_1518 ,           wr_1517 );
  not g2518( wr_1590 ,           wr_1589 );
  not g2519( wr_1700 ,           wr_1699 );
  not g2520( wr_1768 ,           wr_1767 );
  not g2521( G813    ,           wr_1800 );
  nor g2522( wr_2239 , wr_2238 , wr_625  );
  nor g2523( wr_2291 , wr_2290 , wr_625  );
  nor g2524( wr_2569 , wr_2568 , wr_2567 );
  nor g2525( wr_2328 , wr_2327 , wr_2326 );
  nor g2526( wr_2513 , wr_2512 , wr_546  );
  not g2527( wr_2368 ,           wr_2367 );
  nor g2528( wr_2608 , wr_2607 , wr_2606 );
  not g2529( wr_2360 ,           wr_2359 );
  not g2530( wr_2648 ,           wr_2647 );
  not g2531( wr_2640 ,           wr_2639 );
  nor g2532( wr_1371 , wr_1370 , wr_1320 );
  not g2533( wr_1430 ,           wr_1429 );
  nor g2534( wr_1922 , G824    , G4090   );
  nor g2535( wr_1941 , G824    , G4087   );
  nor g2536( wr_1958 , G826    , G4087   );
  nor g2537( wr_1977 , G828    , G4087   );
  nor g2538( wr_1996 , G830    , G4087   );
  nor g2539( wr_2015 , G826    , G4090   );
  nor g2540( wr_2032 , G828    , G4090   );
  nor g2541( wr_2049 , G830    , G4090   );
  nor g2542( wr_2066 , G830    , G1690   );
  nor g2543( wr_2085 , G828    , G1690   );
  nor g2544( wr_2104 , G826    , G1690   );
  nor g2545( wr_2123 , G824    , G1690   );
  nor g2546( wr_2142 , G830    , G1694   );
  nor g2547( wr_2159 , G828    , G1694   );
  nor g2548( wr_2176 , G826    , G1694   );
  nor g2549( wr_2193 , G824    , G1694   );
  not g2550( wr_1486 ,           wr_1485 );
  not g2551( wr_1562 ,           wr_1561 );
  not g2552( wr_1630 ,           wr_1629 );
  not g2553( wr_1706 ,           wr_1705 );
  nor g2554( G863    , wr_1879 , wr_1869 );
  nor g2555( G865    , wr_1892 , wr_1882 );
  nor g2556( G867    , wr_1905 , wr_1895 );
  nor g2557( G869    , wr_1918 , wr_1908 );
  not g2558( wr_1793 ,           wr_1792 );
  not g2559( wr_1483 ,           wr_1482 );
  not g2560( wr_1559 ,           wr_1558 );
  not g2561( wr_1627 ,           wr_1626 );
  not g2562( wr_1703 ,           wr_1702 );
  nor g2563( wr_1519 , wr_1518 , wr_1503 );
  nor g2564( wr_1591 , wr_1590 , wr_1577 );
  nor g2565( wr_1701 , wr_1700 , wr_1685 );
  nor g2566( wr_1769 , wr_1768 , wr_1755 );
  nor g2567( wr_2241 , wr_2240 , wr_2239 );
  nor g2568( wr_2293 , wr_2292 , wr_2291 );
  not g2569( wr_2570 ,           wr_2569 );
  nor g2570( wr_2363 , wr_2328 , wr_2252 );
  nor g2571( wr_2515 , wr_2514 , wr_2513 );
  nor g2572( wr_2572 , wr_2569 , wr_1102 );
  nor g2573( wr_2369 , wr_2368 , wr_2366 );
  nor g2574( wr_2643 , wr_2608 , wr_2526 );
  nor g2575( wr_2329 , wr_2328 , G2174   );
  nor g2576( wr_2361 , wr_2360 , wr_925  );
  nor g2577( wr_2649 , wr_2648 , wr_2646 );
  nor g2578( wr_2609 , wr_2608 , G1497   );
  nor g2579( wr_2641 , wr_2640 , wr_1298 );
  not g2580( wr_1372 ,           wr_1371 );
  nor g2581( wr_1431 , wr_1430 , wr_1392 );
  not g2582( wr_1923 ,           wr_1922 );
  not g2583( wr_1942 ,           wr_1941 );
  not g2584( wr_1959 ,           wr_1958 );
  not g2585( wr_1978 ,           wr_1977 );
  not g2586( wr_1997 ,           wr_1996 );
  not g2587( wr_2016 ,           wr_2015 );
  not g2588( wr_2033 ,           wr_2032 );
  not g2589( wr_2050 ,           wr_2049 );
  not g2590( wr_2067 ,           wr_2066 );
  not g2591( wr_2086 ,           wr_2085 );
  not g2592( wr_2105 ,           wr_2104 );
  not g2593( wr_2124 ,           wr_2123 );
  not g2594( wr_2143 ,           wr_2142 );
  not g2595( wr_2160 ,           wr_2159 );
  not g2596( wr_2177 ,           wr_2176 );
  not g2597( wr_2194 ,           wr_2193 );
  nor g2598( wr_1487 , wr_1486 , G4088   );
  nor g2599( wr_1563 , wr_1562 , G4089   );
  nor g2600( wr_1631 , wr_1630 , G1689   );
  nor g2601( wr_1707 , wr_1706 , G1691   );
  nor g2602( wr_1919 , G863    , G4090   );
  nor g2603( wr_1938 , G863    , G4087   );
  nor g2604( wr_1955 , G865    , G4087   );
  nor g2605( wr_1974 , G867    , G4087   );
  nor g2606( wr_1993 , G869    , G4087   );
  nor g2607( wr_2012 , G865    , G4090   );
  nor g2608( wr_2029 , G867    , G4090   );
  nor g2609( wr_2046 , G869    , G4090   );
  nor g2610( wr_2063 , G869    , G1690   );
  nor g2611( wr_2082 , G867    , G1690   );
  nor g2612( wr_2101 , G865    , G1690   );
  nor g2613( wr_2120 , G863    , G1690   );
  nor g2614( wr_2139 , G869    , G1694   );
  nor g2615( wr_2156 , G867    , G1694   );
  nor g2616( wr_2173 , G865    , G1694   );
  nor g2617( wr_2190 , G863    , G1694   );
  nor g2618( wr_1794 , wr_1793 , wr_1783 );
  nor g2619( wr_1484 , wr_1483 , wr_946  );
  nor g2620( wr_1560 , wr_1559 , wr_1061 );
  nor g2621( wr_1628 , wr_1627 , wr_1442 );
  nor g2622( wr_1704 , wr_1703 , wr_1463 );
  not g2623( G752    ,           wr_1519 );
  not g2624( G792    ,           wr_1591 );
  nor g2625( G670    , wr_1701 , wr_1441 );
  nor g2626( G702    , wr_1769 , wr_1441 );
  not g2627( wr_2242 ,           wr_2241 );
  nor g2628( wr_2244 , wr_2241 , wr_1045 );
  not g2629( wr_2294 ,           wr_2293 );
  nor g2630( wr_2571 , wr_2570 , wr_546  );
  nor g2631( wr_2296 , wr_2293 , wr_1045 );
  not g2632( wr_2364 ,           wr_2363 );
  not g2633( wr_2516 ,           wr_2515 );
  nor g2634( wr_2518 , wr_2515 , wr_1158 );
  not g2635( wr_2644 ,           wr_2643 );
  not g2636( wr_2330 ,           wr_2329 );
  not g2637( wr_2610 ,           wr_2609 );
  nor g2638( wr_1373 , wr_1372 , wr_1306 );
  not g2639( wr_1432 ,           wr_1431 );
  nor g2640( wr_1924 , wr_1923 , G4089   );
  nor g2641( wr_1943 , wr_1942 , G4088   );
  nor g2642( wr_1960 , wr_1959 , G4088   );
  nor g2643( wr_1979 , wr_1978 , G4088   );
  nor g2644( wr_1998 , wr_1997 , G4088   );
  nor g2645( wr_2017 , wr_2016 , G4089   );
  nor g2646( wr_2034 , wr_2033 , G4089   );
  nor g2647( wr_2051 , wr_2050 , G4089   );
  nor g2648( wr_2068 , wr_2067 , G1689   );
  nor g2649( wr_2087 , wr_2086 , G1689   );
  nor g2650( wr_2106 , wr_2105 , G1689   );
  nor g2651( wr_2125 , wr_2124 , G1689   );
  nor g2652( wr_2144 , wr_2143 , G1691   );
  nor g2653( wr_2161 , wr_2160 , G1691   );
  nor g2654( wr_2178 , wr_2177 , G1691   );
  nor g2655( wr_2195 , wr_2194 , G1691   );
  nor g2656( wr_1498 , wr_1497 , wr_1487 );
  nor g2657( wr_1572 , wr_1571 , wr_1563 );
  nor g2658( wr_1642 , wr_1641 , wr_1631 );
  nor g2659( wr_1716 , wr_1715 , wr_1707 );
  not g2660( wr_1920 ,           wr_1919 );
  not g2661( wr_1939 ,           wr_1938 );
  not g2662( wr_1956 ,           wr_1955 );
  not g2663( wr_1975 ,           wr_1974 );
  not g2664( wr_1994 ,           wr_1993 );
  not g2665( wr_2013 ,           wr_2012 );
  not g2666( wr_2030 ,           wr_2029 );
  not g2667( wr_2047 ,           wr_2046 );
  not g2668( wr_2064 ,           wr_2063 );
  not g2669( wr_2083 ,           wr_2082 );
  not g2670( wr_2102 ,           wr_2101 );
  not g2671( wr_2121 ,           wr_2120 );
  not g2672( wr_2140 ,           wr_2139 );
  not g2673( wr_2157 ,           wr_2156 );
  not g2674( wr_2174 ,           wr_2173 );
  not g2675( wr_2191 ,           wr_2190 );
  not g2676( wr_1795 ,           wr_1794 );
  nor g2677( wr_2243 , wr_2242 , wr_610  );
  nor g2678( wr_2295 , wr_2294 , wr_610  );
  nor g2679( wr_2573 , wr_2572 , wr_2571 );
  nor g2680( wr_2365 , wr_2364 , wr_2362 );
  nor g2681( wr_2517 , wr_2516 , wr_538  );
  nor g2682( wr_2645 , wr_2644 , wr_2642 );
  nor g2683( wr_2331 , wr_2330 , wr_854  );
  nor g2684( wr_2611 , wr_2610 , wr_803  );
  not g2685( wr_1374 ,           wr_1373 );
  nor g2686( wr_1433 , wr_1432 , wr_1387 );
  nor g2687( wr_1935 , wr_1934 , wr_1924 );
  nor g2688( wr_1952 , wr_1951 , wr_1943 );
  nor g2689( wr_1971 , wr_1970 , wr_1960 );
  nor g2690( wr_1990 , wr_1989 , wr_1979 );
  nor g2691( wr_2009 , wr_2008 , wr_1998 );
  nor g2692( wr_2026 , wr_2025 , wr_2017 );
  nor g2693( wr_2043 , wr_2042 , wr_2034 );
  nor g2694( wr_2060 , wr_2059 , wr_2051 );
  nor g2695( wr_2079 , wr_2078 , wr_2068 );
  nor g2696( wr_2098 , wr_2097 , wr_2087 );
  nor g2697( wr_2117 , wr_2116 , wr_2106 );
  nor g2698( wr_2136 , wr_2135 , wr_2125 );
  nor g2699( wr_2153 , wr_2152 , wr_2144 );
  nor g2700( wr_2170 , wr_2169 , wr_2161 );
  nor g2701( wr_2187 , wr_2186 , wr_2178 );
  nor g2702( wr_2204 , wr_2203 , wr_2195 );
  not g2703( wr_1499 ,           wr_1498 );
  not g2704( wr_1573 ,           wr_1572 );
  not g2705( wr_1643 ,           wr_1642 );
  not g2706( wr_1717 ,           wr_1716 );
  nor g2707( wr_1921 , wr_1920 , wr_1061 );
  nor g2708( wr_1940 , wr_1939 , wr_946  );
  nor g2709( wr_1957 , wr_1956 , wr_946  );
  nor g2710( wr_1976 , wr_1975 , wr_946  );
  nor g2711( wr_1995 , wr_1994 , wr_946  );
  nor g2712( wr_2014 , wr_2013 , wr_1061 );
  nor g2713( wr_2031 , wr_2030 , wr_1061 );
  nor g2714( wr_2048 , wr_2047 , wr_1061 );
  nor g2715( wr_2065 , wr_2064 , wr_1442 );
  nor g2716( wr_2084 , wr_2083 , wr_1442 );
  nor g2717( wr_2103 , wr_2102 , wr_1442 );
  nor g2718( wr_2122 , wr_2121 , wr_1442 );
  nor g2719( wr_2141 , wr_2140 , wr_1463 );
  nor g2720( wr_2158 , wr_2157 , wr_1463 );
  nor g2721( wr_2175 , wr_2174 , wr_1463 );
  nor g2722( wr_2192 , wr_2191 , wr_1463 );
  nor g2723( wr_1796 , wr_1795 , wr_1780 );
  nor g2724( wr_2245 , wr_2244 , wr_2243 );
  nor g2725( wr_2297 , wr_2296 , wr_2295 );
  not g2726( wr_2574 ,           wr_2573 );
  nor g2727( wr_2370 , wr_2369 , wr_2365 );
  nor g2728( wr_2519 , wr_2518 , wr_2517 );
  nor g2729( wr_2576 , wr_2573 , wr_1158 );
  nor g2730( wr_2650 , wr_2649 , wr_2645 );
  nor g2731( wr_1375 , wr_1374 , wr_1297 );
  not g2732( wr_1434 ,           wr_1433 );
  not g2733( wr_1936 ,           wr_1935 );
  not g2734( wr_1953 ,           wr_1952 );
  not g2735( wr_1972 ,           wr_1971 );
  not g2736( wr_1991 ,           wr_1990 );
  not g2737( wr_2010 ,           wr_2009 );
  not g2738( wr_2027 ,           wr_2026 );
  not g2739( wr_2044 ,           wr_2043 );
  not g2740( wr_2061 ,           wr_2060 );
  not g2741( wr_2080 ,           wr_2079 );
  not g2742( wr_2099 ,           wr_2098 );
  not g2743( wr_2118 ,           wr_2117 );
  not g2744( wr_2137 ,           wr_2136 );
  not g2745( wr_2154 ,           wr_2153 );
  not g2746( wr_2171 ,           wr_2170 );
  not g2747( wr_2188 ,           wr_2187 );
  not g2748( wr_2205 ,           wr_2204 );
  nor g2749( wr_1500 , wr_1499 , wr_1484 );
  nor g2750( wr_1574 , wr_1573 , wr_1560 );
  nor g2751( wr_1644 , wr_1643 , wr_1628 );
  nor g2752( wr_1718 , wr_1717 , wr_1704 );
  nor g2753( G818    , wr_1796 , wr_1772 );
  not g2754( wr_2246 ,           wr_2245 );
  nor g2755( wr_2248 , wr_2245 , wr_1021 );
  not g2756( wr_2298 ,           wr_2297 );
  nor g2757( wr_2575 , wr_2574 , wr_538  );
  nor g2758( wr_2300 , wr_2297 , wr_1021 );
  not g2759( wr_2371 ,           wr_2370 );
  not g2760( wr_2520 ,           wr_2519 );
  nor g2761( wr_2522 , wr_2519 , wr_1134 );
  not g2762( wr_2651 ,           wr_2650 );
  not g2763( wr_1376 ,           wr_1375 );
  nor g2764( wr_1435 , wr_1434 , wr_1386 );
  nor g2765( wr_1937 , wr_1936 , wr_1921 );
  nor g2766( wr_1954 , wr_1953 , wr_1940 );
  nor g2767( wr_1973 , wr_1972 , wr_1957 );
  nor g2768( wr_1992 , wr_1991 , wr_1976 );
  nor g2769( wr_2011 , wr_2010 , wr_1995 );
  nor g2770( wr_2028 , wr_2027 , wr_2014 );
  nor g2771( wr_2045 , wr_2044 , wr_2031 );
  nor g2772( wr_2062 , wr_2061 , wr_2048 );
  nor g2773( wr_2081 , wr_2080 , wr_2065 );
  nor g2774( wr_2100 , wr_2099 , wr_2084 );
  nor g2775( wr_2119 , wr_2118 , wr_2103 );
  nor g2776( wr_2138 , wr_2137 , wr_2122 );
  nor g2777( wr_2155 , wr_2154 , wr_2141 );
  nor g2778( wr_2172 , wr_2171 , wr_2158 );
  nor g2779( wr_2189 , wr_2188 , wr_2175 );
  nor g2780( wr_2206 , wr_2205 , wr_2192 );
  not g2781( G747    ,           wr_1500 );
  not g2782( G787    ,           wr_1574 );
  nor g2783( G642    , wr_1644 , wr_1441 );
  nor g2784( G676    , wr_1718 , wr_1441 );
  nor g2785( wr_2247 , wr_2246 , wr_603  );
  nor g2786( wr_2299 , wr_2298 , wr_603  );
  nor g2787( wr_2577 , wr_2576 , wr_2575 );
  nor g2788( wr_2372 , wr_2371 , wr_2361 );
  nor g2789( wr_2521 , wr_2520 , wr_554  );
  nor g2790( wr_2652 , wr_2651 , wr_2641 );
  nor g2791( wr_1377 , wr_1376 , wr_1296 );
  not g2792( wr_1436 ,           wr_1435 );
  not g2793( G712    ,           wr_1937 );
  not g2794( G727    ,           wr_1954 );
  not g2795( G732    ,           wr_1973 );
  not g2796( G737    ,           wr_1992 );
  not g2797( G742    ,           wr_2011 );
  not g2798( G772    ,           wr_2028 );
  not g2799( G777    ,           wr_2045 );
  not g2800( G782    ,           wr_2062 );
  nor g2801( G645    , wr_2081 , wr_1441 );
  nor g2802( G648    , wr_2100 , wr_1441 );
  nor g2803( G651    , wr_2119 , wr_1441 );
  nor g2804( G654    , wr_2138 , wr_1441 );
  nor g2805( G679    , wr_2155 , wr_1441 );
  nor g2806( G682    , wr_2172 , wr_1441 );
  nor g2807( G685    , wr_2189 , wr_1441 );
  nor g2808( G688    , wr_2206 , wr_1441 );
  nor g2809( wr_2249 , wr_2248 , wr_2247 );
  nor g2810( wr_2301 , wr_2300 , wr_2299 );
  not g2811( wr_2578 ,           wr_2577 );
  not g2812( wr_2373 ,           wr_2372 );
  nor g2813( wr_2523 , wr_2522 , wr_2521 );
  nor g2814( wr_2580 , wr_2577 , wr_1134 );
  not g2815( wr_2653 ,           wr_2652 );
  not g2816( wr_1378 ,           wr_1377 );
  nor g2817( wr_1437 , wr_1436 , wr_1385 );
  not g2818( wr_2250 ,           wr_2249 );
  nor g2819( wr_2302 , wr_2301 , wr_2252 );
  nor g2820( wr_2579 , wr_2578 , wr_554  );
  nor g2821( wr_2374 , wr_2373 , wr_2331 );
  not g2822( wr_2524 ,           wr_2523 );
  nor g2823( wr_2654 , wr_2653 , wr_2611 );
  nor g2824( wr_1379 , wr_1378 , wr_1295 );
  not g2825( wr_1438 ,           wr_1437 );
  nor g2826( wr_2251 , wr_2250 , G2174   );
  nor g2827( wr_2581 , wr_2580 , wr_2579 );
  not g2828( wr_2375 ,           wr_2374 );
  nor g2829( wr_2525 , wr_2524 , G1497   );
  not g2830( wr_2655 ,           wr_2654 );
  not g2831( wr_1380 ,           wr_1379 );
  nor g2832( wr_1439 , wr_1438 , wr_1384 );
  nor g2833( wr_2303 , wr_2302 , wr_2251 );
  nor g2834( wr_2582 , wr_2581 , wr_2526 );
  nor g2835( wr_1381 , wr_1380 , wr_1294 );
  not g2836( wr_1440 ,           wr_1439 );
  not g2837( wr_2377 ,           wr_2303 );
  nor g2838( wr_2376 , wr_2375 , wr_2303 );
  nor g2839( wr_2583 , wr_2582 , wr_2525 );
  not g2840( wr_1382 ,           wr_1381 );
  nor g2841( G585    , wr_1440 , wr_1383 );
  nor g2842( wr_2378 , wr_2374 , wr_2377 );
  not g2843( wr_2657 ,           wr_2583 );
  nor g2844( wr_2656 , wr_2655 , wr_2583 );
  nor g2845( G575    , wr_1382 , wr_1293 );
  nor g2846( wr_2379 , wr_2378 , wr_2376 );
  nor g2847( wr_2658 , wr_2654 , wr_2657 );
  not g2848( wr_2833 ,           wr_2379 );
  nor g2849( wr_2659 , wr_2658 , wr_2656 );
  nor g2850( wr_2380 , wr_2379 , G4092   );
  nor g2851( wr_2834 , wr_2833 , wr_861  );
  not g2852( wr_2822 ,           wr_2659 );
  nor g2853( wr_2660 , wr_2659 , G4092   );
  not g2854( wr_2381 ,           wr_2380 );
  nor g2855( wr_2835 , wr_2834 , wr_2832 );
  nor g2856( wr_2823 , wr_2822 , wr_861  );
  not g2857( wr_2661 ,           wr_2660 );
  nor g2858( wr_2382 , wr_2381 , wr_861  );
  nor g2859( wr_2836 , wr_2835 , G4092   );
  nor g2860( wr_2824 , wr_2823 , wr_2821 );
  nor g2861( wr_2662 , wr_2661 , wr_861  );
  nor g2862( wr_2480 , wr_2479 , wr_2382 );
  nor g2863( wr_2839 , wr_2838 , wr_2836 );
  nor g2864( wr_2825 , wr_2824 , G4092   );
  nor g2865( wr_2820 , wr_2819 , wr_2662 );
  not g2866( G843    ,           wr_2480 );
  nor g2867( wr_2876 , wr_2839 , G1690   );
  nor g2868( wr_2896 , wr_2839 , G1694   );
  nor g2869( wr_2828 , wr_2827 , wr_2825 );
  nor g2870( wr_2840 , wr_2839 , G4087   );
  nor g2871( wr_2859 , wr_2839 , G4090   );
  not g2872( G882    ,           wr_2820 );
  not g2873( wr_2877 ,           wr_2876 );
  not g2874( wr_2897 ,           wr_2896 );
  not g2875( wr_2841 ,           wr_2840 );
  not g2876( wr_2860 ,           wr_2859 );
  nor g2877( wr_2873 , wr_2828 , G1690   );
  nor g2878( wr_2893 , wr_2828 , G1694   );
  nor g2879( wr_2829 , wr_2828 , G4087   );
  nor g2880( wr_2856 , wr_2828 , G4090   );
  nor g2881( wr_2878 , wr_2877 , G1689   );
  nor g2882( wr_2898 , wr_2897 , G1691   );
  nor g2883( wr_2842 , wr_2841 , G4088   );
  nor g2884( wr_2861 , wr_2860 , G4089   );
  not g2885( wr_2874 ,           wr_2873 );
  not g2886( wr_2894 ,           wr_2893 );
  not g2887( wr_2830 ,           wr_2829 );
  not g2888( wr_2857 ,           wr_2856 );
  nor g2889( wr_2889 , wr_2888 , wr_2878 );
  nor g2890( wr_2907 , wr_2906 , wr_2898 );
  nor g2891( wr_2853 , wr_2852 , wr_2842 );
  nor g2892( wr_2870 , wr_2869 , wr_2861 );
  nor g2893( wr_2875 , wr_2874 , wr_1442 );
  nor g2894( wr_2895 , wr_2894 , wr_1463 );
  nor g2895( wr_2831 , wr_2830 , wr_946  );
  nor g2896( wr_2858 , wr_2857 , wr_1061 );
  not g2897( wr_2890 ,           wr_2889 );
  not g2898( wr_2908 ,           wr_2907 );
  not g2899( wr_2854 ,           wr_2853 );
  not g2900( wr_2871 ,           wr_2870 );
  nor g2901( wr_2891 , wr_2890 , wr_2875 );
  nor g2902( wr_2909 , wr_2908 , wr_2895 );
  nor g2903( wr_2855 , wr_2854 , wr_2831 );
  nor g2904( wr_2872 , wr_2871 , wr_2858 );
  nor g2905( wr_2892 , wr_2891 , wr_1441 );
  nor g2906( wr_2910 , wr_2909 , wr_1441 );
  not g2907( G767    ,           wr_2855 );
  not g2908( G807    ,           wr_2872 );
  not g2909( G658    ,           wr_2892 );
  not g2910( G690    ,           wr_2910 );

endmodule
