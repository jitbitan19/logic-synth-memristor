// Benchmark "./input/c3540" written by ABC on Thu Aug  8 02:45:58 2024

module c3540  ( 
    G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116,
    G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200,
    G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274,
    G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698,
    G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107,
    G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190,
    G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270,
    G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_G432_, new_G442_, new_G447_, new_G456_, new_G460_, new_G463_,
    new_G467_, new_G476_, new_G479_, new_G483_, new_G492_, new_G501_,
    new_G504_, new_G513_, new_G517_, new_G526_, new_G530_, new_G540_,
    new_G587_, new_G704_, new_G707_, new_G714_, new_G717_, new_G724_,
    new_G731_, new_G732_, new_G736_, new_G741_, new_G758_, new_G776_,
    new_G780_, new_G788_, new_G791_, new_G798_, new_G799_, new_G802_,
    new_G826_, new_G828_, new_G831_, new_G833_, new_G836_, new_G839_,
    new_G842_, new_G845_, new_G848_, new_G851_, new_G890_, new_G898_,
    new_G907_, new_G1032_, new_G1035_, new_G1048_, new_G1049_, new_G1050_,
    new_G1051_, new_G1540_, new_G1699_, new_G1826_, new_G1827_, new_G1828_,
    new_G2051_, new_G2478_, new_G2865_, new_G2868_, new_G2931_, new_G2934_,
    new_G2939_, new_G2942_, new_G2947_, new_G2950_, new_G2957_, new_G2960_,
    new_G3007_, new_G3079_, new_G3087_, new_G3095_, new_G3103_, new_G3419_,
    new_G588_, new_G759_, new_G1541_, new_G1772_, new_G1829_, new_G1834_,
    new_G2052_, new_G625_, new_G545_, new_G546_, new_G547_, new_G548_,
    new_G549_, new_G550_, new_G551_, new_G552_, new_G2937_, new_G2938_,
    new_G2945_, new_G2946_, new_G621_, new_G626_, new_G635_, new_G636_,
    new_G3085_, new_G3101_, new_G657_, new_G675_, new_G721_, new_G784_,
    new_G794_, new_G807_, new_G816_, new_G823_, new_G860_, new_G861_,
    new_G864_, new_G893_, new_G896_, new_G897_, new_G3093_, new_G905_,
    new_G906_, new_G3109_, new_G973_, new_G980_, new_G987_, new_G994_,
    new_G1001_, new_G1008_, new_G1015_, new_G1022_, new_G1038_, new_G1043_,
    new_G1054_, new_G1057_, new_G1512_, new_G1681_, new_G1717_, new_G1724_,
    new_G1731_, new_G1738_, new_G1745_, new_G1752_, new_G1759_, new_G1766_,
    new_G1773_, new_G1790_, new_G1808_, new_G2278_, new_G2481_, new_G3425_,
    new_G2871_, new_G2874_, new_G2953_, new_G2954_, new_G2963_, new_G2964_,
    new_G3010_, new_G3013_, new_G3017_, new_G3020_, new_G3027_, new_G3030_,
    new_G3037_, new_G3040_, new_G3082_, new_G3090_, new_G3098_, new_G3106_,
    new_G352_, new_G553_, new_G554_, new_G555_, new_G556_, new_G560_,
    new_G561_, new_G650_, new_G956_, new_G974_, new_G975_, new_G976_,
    new_G981_, new_G982_, new_G988_, new_G989_, new_G990_, new_G995_,
    new_G996_, new_G997_, new_G1002_, new_G1003_, new_G1004_, new_G1009_,
    new_G1010_, new_G1016_, new_G1017_, new_G1018_, new_G1023_, new_G1024_,
    new_G1025_, new_G1720_, new_G1727_, new_G1734_, new_G1741_, new_G1748_,
    new_G1755_, new_G1762_, new_G1769_, new_G1791_, new_G1809_, new_G1851_,
    new_G1901_, new_G1952_, new_G2002_, new_G2057_, new_G2109_, new_G2162_,
    new_G2214_, new_G2955_, new_G2956_, new_G2965_, new_G2966_, new_G354_,
    new_G557_, new_G562_, new_G586_, new_G630_, new_G634_, new_G639_,
    new_G642_, new_G3086_, new_G644_, new_G646_, new_G3102_, new_G654_,
    new_G660_, new_G678_, new_G804_, new_G806_, new_G855_, new_G867_,
    new_G903_, new_G3094_, new_G912_, new_G3110_, new_G915_, new_G927_,
    new_G941_, new_G977_, new_G978_, new_G984_, new_G985_, new_G991_,
    new_G992_, new_G998_, new_G999_, new_G1005_, new_G1006_, new_G1012_,
    new_G1013_, new_G1019_, new_G1020_, new_G1026_, new_G1027_, new_G1060_,
    new_G1063_, new_G1066_, new_G1069_, new_G1527_, new_G1530_, new_G1542_,
    new_G1563_, new_G1572_, new_G1581_, new_G1585_, new_G1589_, new_G1593_,
    new_G1597_, new_G1601_, new_G1605_, new_G1716_, new_G1718_, new_G1723_,
    new_G1725_, new_G1730_, new_G1732_, new_G1737_, new_G1739_, new_G1744_,
    new_G1746_, new_G1751_, new_G1753_, new_G1758_, new_G1760_, new_G1765_,
    new_G1767_, new_G1852_, new_G1856_, new_G1870_, new_G1902_, new_G1906_,
    new_G1920_, new_G1953_, new_G1957_, new_G1971_, new_G2003_, new_G2007_,
    new_G2021_, new_G2058_, new_G2062_, new_G2076_, new_G2110_, new_G2114_,
    new_G2128_, new_G2163_, new_G2167_, new_G2181_, new_G2215_, new_G2219_,
    new_G2233_, new_G2285_, new_G2288_, new_G2289_, new_G2293_, new_G2298_,
    new_G2302_, new_G2877_, new_G2983_, new_G2986_, new_G3014_, new_G3015_,
    new_G3023_, new_G3024_, new_G3033_, new_G3034_, new_G3043_, new_G3044_,
    new_G643_, new_G647_, new_G680_, new_G904_, new_G913_, new_G920_,
    new_G979_, new_G993_, new_G1000_, new_G1007_, new_G1021_, new_G1028_,
    new_G1719_, new_G1721_, new_G1726_, new_G1728_, new_G1733_, new_G1735_,
    new_G1740_, new_G1742_, new_G1747_, new_G1749_, new_G1754_, new_G1756_,
    new_G1761_, new_G1763_, new_G1768_, new_G1770_, new_G1794_, new_G1799_,
    new_G1812_, new_G1817_, new_G1859_, new_G1909_, new_G1960_, new_G2010_,
    new_G2065_, new_G2117_, new_G2170_, new_G2222_, new_G2678_, new_G2697_,
    new_G2716_, new_G2733_, new_G2751_, new_G2768_, new_G2785_, new_G2802_,
    new_G3016_, new_G3025_, new_G3026_, new_G3035_, new_G3036_, new_G3045_,
    new_G3046_, new_G2989_, new_G2990_, new_G610_, new_G613_, new_G616_,
    new_G640_, new_G648_, new_G655_, new_G665_, new_G668_, new_G671_,
    new_G683_, new_G685_, new_G688_, new_G694_, new_G696_, new_G699_,
    new_G870_, new_G887_, new_G901_, new_G910_, new_G914_, new_G916_,
    new_G942_, new_G943_, new_G1072_, new_G1084_, new_G1096_, new_G1108_,
    new_G1120_, new_G1132_, new_G1144_, new_G1156_, new_G1533_, new_G1534_,
    new_G1535_, new_G1545_, new_G1554_, new_G1610_, new_G1619_, new_G1628_,
    new_G1637_, new_G1646_, new_G1655_, new_G1664_, new_G1673_, new_G1722_,
    new_G1729_, new_G1736_, new_G1743_, new_G1750_, new_G1757_, new_G1764_,
    new_G1771_, new_G1853_, new_G1954_, new_G2004_, new_G2059_, new_G2164_,
    new_G2216_, new_G2485_, new_G2900_, new_G2903_, new_G2967_, new_G2970_,
    new_G2975_, new_G2978_, new_G3047_, new_G3050_, new_G3055_, new_G3058_,
    new_G574_, new_G575_, new_G617_, new_G641_, new_G649_, new_G662_,
    new_G672_, new_G690_, new_G691_, new_G701_, new_G702_, new_G902_,
    new_G911_, new_G917_, new_G923_, new_G1538_, new_G1871_, new_G1872_,
    new_G1873_, new_G1921_, new_G1922_, new_G1923_, new_G1972_, new_G1973_,
    new_G1974_, new_G2022_, new_G2023_, new_G2024_, new_G2077_, new_G2078_,
    new_G2079_, new_G2129_, new_G2130_, new_G2131_, new_G2182_, new_G2183_,
    new_G2184_, new_G2234_, new_G2235_, new_G2236_, new_G2973_, new_G2974_,
    new_G2981_, new_G2982_, new_G576_, new_G3053_, new_G3054_, new_G3061_,
    new_G3062_, new_G645_, new_G926_, new_G928_, new_G947_, new_G983_,
    new_G1011_, new_G1075_, new_G1087_, new_G1099_, new_G1111_, new_G1123_,
    new_G1135_, new_G1147_, new_G1159_, new_G1168_, new_G1177_, new_G1186_,
    new_G1195_, new_G1204_, new_G1213_, new_G1222_, new_G1231_, new_G1609_,
    new_G1611_, new_G1618_, new_G1620_, new_G1627_, new_G1629_, new_G1636_,
    new_G1638_, new_G1645_, new_G1647_, new_G1654_, new_G1656_, new_G1663_,
    new_G1665_, new_G1672_, new_G1674_, new_G1862_, new_G1866_, new_G1874_,
    new_G1924_, new_G1963_, new_G1967_, new_G1975_, new_G2013_, new_G2017_,
    new_G2025_, new_G2068_, new_G2072_, new_G2080_, new_G2132_, new_G2173_,
    new_G2177_, new_G2185_, new_G2225_, new_G2229_, new_G2237_, new_G2488_,
    new_G2679_, new_G2680_, new_G2698_, new_G2699_, new_G2717_, new_G2718_,
    new_G2734_, new_G2735_, new_G2752_, new_G2753_, new_G2769_, new_G2770_,
    new_G2786_, new_G2787_, new_G2803_, new_G2804_, new_G359_, new_G1029_,
    new_G565_, new_G566_, new_G569_, new_G570_, new_G589_, new_G590_,
    new_G595_, new_G596_, new_G929_, new_G938_, new_G944_, new_G986_,
    new_G1014_, new_G1616_, new_G1625_, new_G1634_, new_G1643_, new_G360_,
    new_G567_, new_G571_, new_G579_, new_G591_, new_G597_, new_G614_,
    new_G1240_, new_G1241_, new_G1242_, new_G1243_, new_G1244_, new_G1245_,
    new_G1246_, new_G1247_, new_G1257_, new_G1258_, new_G1259_, new_G1260_,
    new_G1261_, new_G1262_, new_G1263_, new_G1264_, new_G1274_, new_G1275_,
    new_G1276_, new_G1277_, new_G1278_, new_G1279_, new_G1280_, new_G1281_,
    new_G1291_, new_G1292_, new_G1293_, new_G1294_, new_G1295_, new_G1296_,
    new_G1297_, new_G1298_, new_G1308_, new_G1309_, new_G1310_, new_G1311_,
    new_G1312_, new_G1313_, new_G1314_, new_G1315_, new_G1325_, new_G1326_,
    new_G1327_, new_G1328_, new_G1329_, new_G1330_, new_G1331_, new_G1332_,
    new_G1342_, new_G1343_, new_G1344_, new_G1345_, new_G1346_, new_G1347_,
    new_G1348_, new_G1349_, new_G1359_, new_G1360_, new_G1361_, new_G1362_,
    new_G1363_, new_G1364_, new_G1365_, new_G1366_, new_G1376_, new_G1377_,
    new_G1378_, new_G1379_, new_G1380_, new_G1381_, new_G1382_, new_G1383_,
    new_G1393_, new_G1394_, new_G1395_, new_G1396_, new_G1397_, new_G1398_,
    new_G1399_, new_G1400_, new_G1410_, new_G1411_, new_G1412_, new_G1413_,
    new_G1414_, new_G1415_, new_G1416_, new_G1417_, new_G1427_, new_G1428_,
    new_G1429_, new_G1430_, new_G1431_, new_G1432_, new_G1433_, new_G1434_,
    new_G1444_, new_G1445_, new_G1446_, new_G1447_, new_G1448_, new_G1449_,
    new_G1450_, new_G1451_, new_G1461_, new_G1462_, new_G1463_, new_G1464_,
    new_G1465_, new_G1466_, new_G1467_, new_G1468_, new_G1478_, new_G1479_,
    new_G1480_, new_G1481_, new_G1482_, new_G1483_, new_G1484_, new_G1485_,
    new_G1495_, new_G1496_, new_G1497_, new_G1498_, new_G1499_, new_G1500_,
    new_G1501_, new_G1502_, new_G1877_, new_G1880_, new_G1891_, new_G1903_,
    new_G1927_, new_G1930_, new_G1978_, new_G1981_, new_G1992_, new_G2028_,
    new_G2031_, new_G2042_, new_G2085_, new_G2088_, new_G2099_, new_G2111_,
    new_G2137_, new_G2140_, new_G2190_, new_G2193_, new_G2204_, new_G2242_,
    new_G2245_, new_G2256_, new_G2320_, new_G2341_, new_G2354_, new_G2367_,
    new_G2383_, new_G2391_, new_G2474_, new_G2475_, new_G2476_, new_G2477_,
    new_G2482_, new_G568_, new_G618_, new_G1248_, new_G1249_, new_G1250_,
    new_G1251_, new_G1252_, new_G1253_, new_G1254_, new_G1255_, new_G1265_,
    new_G1266_, new_G1267_, new_G1268_, new_G1269_, new_G1270_, new_G1271_,
    new_G1272_, new_G1282_, new_G1283_, new_G1284_, new_G1285_, new_G1286_,
    new_G1287_, new_G1288_, new_G1289_, new_G1299_, new_G1300_, new_G1301_,
    new_G1302_, new_G1303_, new_G1304_, new_G1305_, new_G1306_, new_G1316_,
    new_G1317_, new_G1318_, new_G1319_, new_G1320_, new_G1321_, new_G1322_,
    new_G1323_, new_G1333_, new_G1334_, new_G1335_, new_G1336_, new_G1337_,
    new_G1338_, new_G1339_, new_G1340_, new_G1350_, new_G1351_, new_G1352_,
    new_G1353_, new_G1354_, new_G1355_, new_G1356_, new_G1357_, new_G1367_,
    new_G1368_, new_G1369_, new_G1370_, new_G1371_, new_G1372_, new_G1373_,
    new_G1374_, new_G1384_, new_G1385_, new_G1386_, new_G1387_, new_G1388_,
    new_G1389_, new_G1390_, new_G1391_, new_G1401_, new_G1402_, new_G1403_,
    new_G1404_, new_G1405_, new_G1406_, new_G1407_, new_G1408_, new_G1418_,
    new_G1419_, new_G1420_, new_G1421_, new_G1422_, new_G1423_, new_G1424_,
    new_G1425_, new_G1435_, new_G1436_, new_G1437_, new_G1438_, new_G1439_,
    new_G1440_, new_G1441_, new_G1442_, new_G1452_, new_G1453_, new_G1454_,
    new_G1455_, new_G1456_, new_G1457_, new_G1458_, new_G1459_, new_G1469_,
    new_G1470_, new_G1471_, new_G1472_, new_G1473_, new_G1474_, new_G1475_,
    new_G1476_, new_G1486_, new_G1487_, new_G1488_, new_G1489_, new_G1490_,
    new_G1491_, new_G1492_, new_G1493_, new_G1503_, new_G1504_, new_G1505_,
    new_G1506_, new_G1507_, new_G1508_, new_G1509_, new_G1510_, new_G2483_,
    new_G600_, new_G661_, new_G669_, new_G679_, new_G1256_, new_G1273_,
    new_G1290_, new_G1307_, new_G1324_, new_G1341_, new_G1358_, new_G1375_,
    new_G1392_, new_G1409_, new_G1426_, new_G1443_, new_G1460_, new_G1477_,
    new_G1494_, new_G1511_, new_G1652_, new_G1883_, new_G1886_, new_G1889_,
    new_G1890_, new_G1912_, new_G1916_, new_G1984_, new_G1987_, new_G1990_,
    new_G1991_, new_G2034_, new_G2037_, new_G2040_, new_G2041_, new_G2091_,
    new_G2094_, new_G2097_, new_G2098_, new_G2120_, new_G2124_, new_G2196_,
    new_G2199_, new_G2202_, new_G2203_, new_G2248_, new_G2251_, new_G2254_,
    new_G2255_, new_G2484_, new_G2991_, new_G2994_, new_G2999_, new_G3002_,
    new_G3063_, new_G3071_, new_G3124_, new_G3134_, new_G3158_, new_G3166_,
    new_G3174_, new_G3182_, new_G3190_, new_G3200_, new_G3224_, new_G3232_,
    new_G3240_, new_G3248_, new_G663_, new_G673_, new_G681_, new_G1536_,
    new_G1537_, new_G1582_, new_G1583_, new_G1586_, new_G1587_, new_G1590_,
    new_G1591_, new_G1594_, new_G1595_, new_G1598_, new_G1599_, new_G1602_,
    new_G1603_, new_G1606_, new_G1607_, new_G1894_, new_G1997_, new_G2047_,
    new_G2102_, new_G2209_, new_G2261_, new_G2489_, new_G3005_, new_G3006_,
    new_G3077_, new_G3069_, new_G2997_, new_G2998_, new_G689_, new_G700_,
    new_G1539_, new_G1584_, new_G1588_, new_G1592_, new_G1596_, new_G1600_,
    new_G1604_, new_G1608_, new_G1661_, new_G1892_, new_G1893_, new_G1933_,
    new_G1936_, new_G1939_, new_G1940_, new_G1941_, new_G1993_, new_G1996_,
    new_G2043_, new_G2046_, new_G2100_, new_G2101_, new_G2143_, new_G2146_,
    new_G2149_, new_G2150_, new_G2151_, new_G2205_, new_G2208_, new_G2257_,
    new_G2260_, new_G3138_, new_G2328_, new_G3162_, new_G3170_, new_G3178_,
    new_G3186_, new_G3204_, new_G2375_, new_G3236_, new_G3244_, new_G3252_,
    new_G3228_, new_G3066_, new_G3074_, new_G3128_, new_G3194_, new_G619_,
    new_G620_, new_G582_, new_G583_, new_G692_, new_G703_, new_G1612_,
    new_G1621_, new_G1630_, new_G1639_, new_G1648_, new_G1657_, new_G1666_,
    new_G1675_, new_G1895_, new_G1946_, new_G1998_, new_G2048_, new_G2103_,
    new_G2156_, new_G2210_, new_G2262_, new_G2271_, new_G2311_, new_G356_,
    new_G357_, new_G603_, new_G3078_, new_G606_, new_G3070_, new_G1670_,
    new_G1679_, new_G1942_, new_G1945_, new_G2152_, new_G2155_, new_G2445_,
    new_G2448_, new_G2455_, new_G2458_, new_G3142_, new_G3150_, new_G3208_,
    new_G3216_, new_G604_, new_G607_, new_G1947_, new_G2157_, new_G2317_,
    new_G2338_, new_G2351_, new_G2364_, new_G2380_, new_G2388_, new_G605_,
    new_G608_, new_G2272_, new_G2312_, new_G3146_, new_G3154_, new_G3220_,
    new_G3212_, new_G2444_, new_G2451_, new_G2454_, new_G2461_, new_G2530_,
    new_G3323_, new_G349_, new_G350_, new_G2265_, new_G2273_, new_G2274_,
    new_G2309_, new_G2313_, new_G2314_, new_G2325_, new_G2372_, new_G2523_,
    new_G2533_, new_G3121_, new_G3131_, new_G3155_, new_G3163_, new_G3171_,
    new_G3179_, new_G3187_, new_G3197_, new_G3221_, new_G3229_, new_G3237_,
    new_G3245_, new_G2275_, new_G2315_, new_G3329_, new_G2324_, new_G2350_,
    new_G2363_, new_G2371_, new_G2387_, new_G2400_, new_G2268_, new_G3137_,
    new_G3161_, new_G2345_, new_G3169_, new_G3177_, new_G2358_, new_G3185_,
    new_G3203_, new_G3235_, new_G3243_, new_G2395_, new_G3251_, new_G3227_,
    new_G2432_, new_G2490_, new_G3127_, new_G3130_, new_G3139_, new_G3147_,
    new_G3193_, new_G3196_, new_G3205_, new_G3213_, new_G2307_, new_G2308_,
    new_G2323_, new_G2349_, new_G2362_, new_G2370_, new_G2386_, new_G2399_,
    new_G2344_, new_G2357_, new_G2394_, new_G2431_, new_G2464_, new_G2491_,
    new_G3129_, new_G3195_, new_G368_, new_G1615_, new_G2337_, new_G1633_,
    new_G1642_, new_G1651_, new_G2379_, new_G1669_, new_G1678_, new_G3145_,
    new_G2332_, new_G3153_, new_G2346_, new_G2359_, new_G3219_, new_G2396_,
    new_G3211_, new_G2425_, new_G2433_, new_G3272_, new_G3308_, new_G1613_,
    new_G2336_, new_G1631_, new_G1640_, new_G1649_, new_G2378_, new_G1667_,
    new_G1676_, new_G2331_, new_G2424_, new_G2467_, new_G2495_, new_G3295_,
    new_G3374_, new_G1614_, new_G1624_, new_G1632_, new_G1641_, new_G1650_,
    new_G1660_, new_G1668_, new_G1677_, new_G2333_, new_G2406_, new_G2409_,
    new_G2415_, new_G2419_, new_G2426_, new_G2439_, new_G2518_, new_G3276_,
    new_G3312_, new_G2612_, new_G3326_, new_G1617_, new_G1622_, new_G1635_,
    new_G1644_, new_G1653_, new_G1658_, new_G1671_, new_G1680_, new_G2500_,
    new_G2505_, new_G2519_, new_G3378_, new_G2642_, new_G2645_, new_G3301_,
    new_G1623_, new_G1659_, new_G2401_, new_G2501_, new_G2511_, new_G2512_,
    new_G2513_, new_G2514_, new_G2517_, new_G2531_, new_G2532_, new_G2534_,
    new_G2535_, new_G2607_, new_G3330_, new_G2643_, new_G2687_, new_G2725_,
    new_G2742_, new_G2760_, new_G2794_, new_G2811_, new_G3280_, new_G3290_,
    new_G3298_, new_G3316_, new_G3406_, new_G3414_, new_G3422_, new_G1626_,
    new_G1662_, new_G2567_, new_G2589_, new_G2608_, new_G2654_, new_G3253_,
    new_G3277_, new_G3287_, new_G3305_, new_G3313_, new_G3350_, new_G932_,
    new_G2508_, new_G2524_, new_G2525_, new_G2526_, new_G3294_, new_G2609_,
    new_G3410_, new_G3418_, new_G2624_, new_G3426_, new_G2629_, new_G2647_,
    new_G2706_, new_G2777_, new_G3264_, new_G3284_, new_G3302_, new_G3303_,
    new_G3320_, new_G3398_, new_G2657_, new_G398_, new_G933_, new_G2527_,
    new_G3259_, new_G3354_, new_G3293_, new_G2563_, new_G3311_, new_G2585_,
    new_G2625_, new_G3283_, new_G3286_, new_G3304_, new_G3319_, new_G3322_,
    new_G3358_, new_G3366_, new_G3382_, new_G3390_, new_G397_, new_G2544_,
    new_G2562_, new_G2584_, new_G3402_, new_G2626_, new_G2632_, new_G2634_,
    new_G2650_, new_G3268_, new_G3256_, new_G3285_, new_G3321_, new_G3371_,
    new_G3403_, new_G3411_, new_G362_, new_G1030_, new_G2564_, new_G3362_,
    new_G3370_, new_G2586_, new_G3386_, new_G3394_, new_G2633_, new_G3261_,
    new_G3269_, new_G3347_, new_G3395_, new_G363_, new_G2536_, new_G3260_,
    new_G3377_, new_G2580_, new_G3409_, new_G2616_, new_G3417_, new_G2622_,
    new_G2635_, new_G2805_, new_G2808_, new_G3334_, new_G3342_, new_G3454_,
    new_G2537_, new_G3275_, new_G2540_, new_G3353_, new_G2557_, new_G2579_,
    new_G3401_, new_G2602_, new_G2615_, new_G2621_, new_G3267_, new_G3112_,
    new_G3355_, new_G3363_, new_G3379_, new_G3387_, new_G2538_, new_G2539_,
    new_G3338_, new_G3346_, new_G2556_, new_G2581_, new_G2601_, new_G2617_,
    new_G2623_, new_G2638_, new_G3458_, new_G2814_, new_G2816_, new_G3111_,
    new_G2541_, new_G2558_, new_G3361_, new_G2571_, new_G3369_, new_G2577_,
    new_G3385_, new_G2593_, new_G3393_, new_G2598_, new_G2603_, new_G3113_,
    new_G3116_, new_G3451_, new_G395_, new_G2570_, new_G2576_, new_G2592_,
    new_G2597_, new_G2736_, new_G2739_, new_G2788_, new_G3438_, new_G3446_,
    new_G3459_, new_G3119_, new_G3120_, new_G2572_, new_G2578_, new_G2594_,
    new_G2599_, new_G2677_, new_G3457_, new_G2700_, new_G2771_, new_G3331_,
    new_G3339_, new_G3427_, new_G3443_, new_G954_, new_G955_, new_G2600_,
    new_G3442_, new_G3450_, new_G2676_, new_G2745_, new_G2748_, new_G3465_,
    new_G3435_, new_G950_, new_G3337_, new_G2548_, new_G3345_, new_G2553_,
    new_G2661_, new_G2662_, new_G3433_, new_G3449_, new_G2672_, new_G2674_,
    new_G2719_, new_G2754_, new_G3430_, new_G383_, new_G951_, new_G2547_,
    new_G2552_, new_G2663_, new_G2670_, new_G3441_, new_G2671_, new_G2675_,
    new_G3491_, new_G3499_, new_G2549_, new_G2554_, new_G2664_, new_G3434_,
    new_G2669_, new_G2673_, new_G2757_, new_G2791_, new_G365_, new_G1031_,
    new_G2555_, new_G2665_, new_G2667_, new_G2774_, new_G3497_, new_G3505_,
    new_G366_, new_G2658_, new_G2659_, new_G2666_, new_G2668_, new_G2681_,
    new_G2763_, new_G2765_, new_G2797_, new_G2799_, new_G2660_, new_G2703_,
    new_G2722_, new_G2780_, new_G2782_, new_G386_, new_G392_, new_G2684_,
    new_G3462_, new_G3470_, new_G389_, new_G2709_, new_G2713_, new_G2728_,
    new_G2730_, new_G2922_, new_G3467_, new_G2690_, new_G2694_, new_G2821_,
    new_G3466_, new_G3474_, new_G380_, new_G2822_, new_G3473_, new_G2827_,
    new_G2839_, new_G2883_, new_G3507_, new_G2823_, new_G2826_, new_G2880_,
    new_G2925_, new_G2928_, new_G3510_, new_G2828_, new_G3494_, new_G3502_,
    new_G3513_, new_G3544_, new_G3552_, new_G406_, new_G2929_, new_G3475_,
    new_G3483_, new_G3514_, new_G3515_, new_G3541_, new_G3549_, new_G2930_,
    new_G2842_, new_G3498_, new_G2852_, new_G3506_, new_G3548_, new_G3556_,
    new_G3478_, new_G3486_, new_G3516_, new_G408_, new_G3481_, new_G3489_,
    new_G2843_, new_G2853_, new_G3547_, new_G2887_, new_G2896_, new_G3555_,
    new_G3520_, new_G2831_, new_G3482_, new_G2836_, new_G3490_, new_G2844_,
    new_G2848_, new_G2886_, new_G2895_, new_G2832_, new_G2837_, new_G2849_,
    new_G3524_, new_G2888_, new_G2891_, new_G2833_, new_G2838_, new_G2892_,
    new_G3517_, new_G2906_, new_G2908_, new_G2913_, new_G3523_, new_G2855_,
    new_G2907_, new_G2909_, new_G3525_, new_G3533_, new_G2854_, new_G2910_,
    new_G3560_, new_G3568_, new_G2856_, new_G3539_, new_G3531_, new_G3572_,
    new_G3564_, new_G3557_, new_G3565_, new_G3528_, new_G3536_, new_G2921_,
    new_G2917_, new_G3571_, new_G3563_, new_G2863_, new_G2859_, new_G2920_,
    new_G2916_, new_G3540_, new_G3532_, new_G2864_, new_G2860_, new_G403_,
    new_G404_, new_G400_, new_G401_;
  assign new_G432_ = G50;
  assign new_G442_ = ~G50;
  assign new_G447_ = G58;
  assign new_G456_ = ~G58;
  assign new_G460_ = G68;
  assign new_G463_ = ~G68;
  assign new_G467_ = G68;
  assign new_G476_ = G77;
  assign new_G479_ = ~G77;
  assign new_G483_ = G77;
  assign new_G492_ = G87;
  assign new_G501_ = ~G87;
  assign new_G504_ = G97;
  assign new_G513_ = ~G97;
  assign new_G517_ = G107;
  assign new_G526_ = ~G107;
  assign new_G530_ = G116;
  assign new_G540_ = ~G116;
  assign new_G587_ = G257 | G264;
  assign new_G704_ = ~G1;
  assign new_G707_ = G1;
  assign new_G714_ = ~G1;
  assign new_G717_ = G13;
  assign new_G724_ = ~G13;
  assign new_G731_ = G13 & G20;
  assign new_G732_ = ~G20;
  assign new_G736_ = G20;
  assign new_G741_ = ~G20;
  assign new_G758_ = ~G33;
  assign new_G776_ = G33;
  assign new_G780_ = ~G33;
  assign new_G788_ = G33 & G41;
  assign new_G791_ = ~G41;
  assign new_G798_ = G41 | G45;
  assign new_G799_ = G45;
  assign new_G802_ = ~G45;
  assign new_G826_ = ~G50;
  assign new_G828_ = G58;
  assign new_G831_ = ~G58;
  assign new_G833_ = G68;
  assign new_G836_ = ~G68;
  assign new_G839_ = G87;
  assign new_G842_ = ~G87;
  assign new_G845_ = G97;
  assign new_G848_ = ~G97;
  assign new_G851_ = ~G107;
  assign new_G890_ = G1;
  assign new_G898_ = G68;
  assign new_G907_ = G107;
  assign new_G1032_ = ~G20;
  assign new_G1035_ = G190;
  assign new_G1048_ = ~G200;
  assign new_G1049_ = G20 & G200;
  assign new_G1050_ = ~G20 | ~G200;
  assign new_G1051_ = G20 & G179;
  assign new_G1540_ = ~G20;
  assign new_G1699_ = G1698 | G33;
  assign new_G1826_ = ~G1 | ~G13;
  assign new_G1827_ = ~G33 | ~G1 | ~G20;
  assign new_G1828_ = ~G20;
  assign new_G2051_ = ~G33;
  assign new_G2478_ = G179;
  assign new_G2865_ = ~G213;
  assign new_G2868_ = G343;
  assign new_G2931_ = G226;
  assign new_G2934_ = G232;
  assign new_G2939_ = G238;
  assign new_G2942_ = G244;
  assign new_G2947_ = G250;
  assign new_G2950_ = G257;
  assign new_G2957_ = G264;
  assign new_G2960_ = G270;
  assign new_G3007_ = G50;
  assign new_G3079_ = G58;
  assign new_G3087_ = G58;
  assign new_G3095_ = G97;
  assign new_G3103_ = G97;
  assign new_G3419_ = G330;
  assign new_G588_ = G250 & new_G587_;
  assign new_G759_ = new_G758_ | G20;
  assign new_G1541_ = new_G1540_ | G169;
  assign new_G1772_ = ~new_G731_;
  assign new_G1829_ = new_G1828_ | G1;
  assign new_G1834_ = new_G1826_ & new_G1827_;
  assign new_G2052_ = new_G2051_ | G1;
  assign new_G625_ = new_G836_ & new_G826_ & new_G831_;
  assign new_G545_ = ~G226 | ~new_G432_;
  assign new_G546_ = ~G232 | ~new_G447_;
  assign new_G547_ = ~G238 | ~new_G467_;
  assign new_G548_ = ~G244 | ~new_G483_;
  assign new_G549_ = ~G250 | ~new_G492_;
  assign new_G550_ = ~G257 | ~new_G504_;
  assign new_G551_ = ~G264 | ~new_G517_;
  assign new_G552_ = ~G270 | ~new_G530_;
  assign new_G2937_ = ~new_G2931_;
  assign new_G2938_ = ~new_G2934_;
  assign new_G2945_ = ~new_G2939_;
  assign new_G2946_ = ~new_G2942_;
  assign new_G621_ = ~new_G456_ | ~new_G463_;
  assign new_G626_ = ~new_G513_ | ~new_G526_;
  assign new_G635_ = ~new_G460_ | ~new_G476_;
  assign new_G636_ = new_G442_;
  assign new_G3085_ = ~new_G3079_;
  assign new_G3101_ = ~new_G3095_;
  assign new_G657_ = new_G802_;
  assign new_G675_ = new_G802_;
  assign new_G721_ = new_G717_;
  assign new_G784_ = new_G780_;
  assign new_G794_ = new_G791_;
  assign new_G807_ = new_G714_ & new_G798_;
  assign new_G816_ = new_G791_ & new_G714_ & new_G799_;
  assign new_G823_ = new_G704_ & new_G799_;
  assign new_G860_ = new_G736_ & new_G707_ & new_G724_;
  assign new_G861_ = ~new_G736_ | ~new_G707_ | ~new_G724_;
  assign new_G864_ = ~new_G707_ | ~new_G724_;
  assign new_G893_ = new_G890_;
  assign new_G896_ = ~G45 | ~new_G717_ | ~new_G732_;
  assign new_G897_ = ~new_G836_ | ~new_G826_ | ~new_G831_;
  assign new_G3093_ = ~new_G3087_;
  assign new_G905_ = new_G851_ & new_G842_ & new_G848_;
  assign new_G906_ = ~new_G851_ | ~new_G842_ | ~new_G848_;
  assign new_G3109_ = ~new_G3103_;
  assign new_G973_ = ~new_G741_;
  assign new_G980_ = ~new_G741_;
  assign new_G987_ = ~new_G741_;
  assign new_G994_ = ~new_G741_;
  assign new_G1001_ = ~new_G741_;
  assign new_G1008_ = ~new_G741_;
  assign new_G1015_ = ~new_G741_;
  assign new_G1022_ = ~new_G741_;
  assign new_G1038_ = new_G1032_ | new_G1035_;
  assign new_G1043_ = ~new_G1032_ & ~new_G1035_;
  assign new_G1054_ = new_G1051_;
  assign new_G1057_ = ~new_G1051_;
  assign new_G1512_ = new_G776_;
  assign new_G1681_ = new_G780_;
  assign new_G1717_ = ~new_G1699_;
  assign new_G1724_ = ~new_G1699_;
  assign new_G1731_ = ~new_G1699_;
  assign new_G1738_ = ~new_G1699_;
  assign new_G1745_ = ~new_G1699_;
  assign new_G1752_ = ~new_G1699_;
  assign new_G1759_ = ~new_G1699_;
  assign new_G1766_ = ~new_G1699_;
  assign new_G1773_ = G1 | new_G1772_;
  assign new_G1790_ = ~new_G788_;
  assign new_G1808_ = ~new_G788_;
  assign new_G2278_ = new_G732_ & new_G704_ & new_G717_;
  assign new_G2481_ = ~new_G2478_;
  assign new_G3425_ = ~new_G3419_;
  assign new_G2871_ = new_G2865_ | new_G2868_;
  assign new_G2874_ = ~new_G2865_ & ~new_G2868_;
  assign new_G2953_ = ~new_G2947_;
  assign new_G2954_ = ~new_G2950_;
  assign new_G2963_ = ~new_G2957_;
  assign new_G2964_ = ~new_G2960_;
  assign new_G3010_ = new_G456_;
  assign new_G3013_ = ~new_G3007_;
  assign new_G3017_ = new_G463_;
  assign new_G3020_ = new_G479_;
  assign new_G3027_ = new_G501_;
  assign new_G3030_ = new_G513_;
  assign new_G3037_ = new_G526_;
  assign new_G3040_ = new_G540_;
  assign new_G3082_ = new_G898_;
  assign new_G3090_ = new_G898_;
  assign new_G3098_ = new_G907_;
  assign new_G3106_ = new_G907_;
  assign new_G352_ = ~new_G479_ | ~new_G625_;
  assign new_G553_ = new_G548_ & new_G547_ & new_G545_ & new_G546_;
  assign new_G554_ = new_G552_ & new_G551_ & new_G549_ & new_G550_;
  assign new_G555_ = ~new_G2934_ | ~new_G2937_;
  assign new_G556_ = ~new_G2931_ | ~new_G2938_;
  assign new_G560_ = ~new_G2942_ | ~new_G2945_;
  assign new_G561_ = ~new_G2939_ | ~new_G2946_;
  assign new_G650_ = new_G432_ & new_G621_;
  assign new_G956_ = new_G890_ & new_G896_;
  assign new_G974_ = ~new_G759_;
  assign new_G975_ = new_G741_ & new_G759_;
  assign new_G976_ = new_G897_ & new_G973_;
  assign new_G981_ = ~new_G759_;
  assign new_G982_ = new_G741_ & new_G759_;
  assign new_G988_ = ~new_G759_;
  assign new_G989_ = new_G741_ & new_G759_;
  assign new_G990_ = new_G836_ & new_G987_;
  assign new_G995_ = ~new_G759_;
  assign new_G996_ = new_G741_ & new_G759_;
  assign new_G997_ = G77 & new_G994_;
  assign new_G1002_ = ~new_G759_;
  assign new_G1003_ = new_G741_ & new_G759_;
  assign new_G1004_ = new_G906_ & new_G1001_;
  assign new_G1009_ = ~new_G759_;
  assign new_G1010_ = new_G741_ & new_G759_;
  assign new_G1016_ = ~new_G759_;
  assign new_G1017_ = new_G741_ & new_G759_;
  assign new_G1018_ = new_G851_ & new_G1015_;
  assign new_G1023_ = ~new_G759_;
  assign new_G1024_ = new_G741_ & new_G759_;
  assign new_G1025_ = G116 & new_G1022_;
  assign new_G1720_ = G222 & new_G1717_;
  assign new_G1727_ = G223 & new_G1724_;
  assign new_G1734_ = G226 & new_G1731_;
  assign new_G1741_ = G232 & new_G1738_;
  assign new_G1748_ = G238 & new_G1745_;
  assign new_G1755_ = G244 & new_G1752_;
  assign new_G1762_ = G250 & new_G1759_;
  assign new_G1769_ = G257 & new_G1766_;
  assign new_G1791_ = new_G1790_ & G1 & G13;
  assign new_G1809_ = new_G1808_ & G1 & G13;
  assign new_G1851_ = ~new_G1834_;
  assign new_G1901_ = ~new_G1834_;
  assign new_G1952_ = ~new_G1834_;
  assign new_G2002_ = ~new_G1834_;
  assign new_G2057_ = ~new_G1834_;
  assign new_G2109_ = ~new_G1834_;
  assign new_G2162_ = ~new_G1834_;
  assign new_G2214_ = ~new_G1834_;
  assign new_G2955_ = ~new_G2950_ | ~new_G2953_;
  assign new_G2956_ = ~new_G2947_ | ~new_G2954_;
  assign new_G2965_ = ~new_G2960_ | ~new_G2963_;
  assign new_G2966_ = ~new_G2957_ | ~new_G2964_;
  assign G353 = ~new_G352_;
  assign new_G354_ = G87 & new_G626_;
  assign new_G557_ = ~new_G555_ | ~new_G556_;
  assign new_G562_ = ~new_G560_ | ~new_G561_;
  assign new_G586_ = ~new_G553_ | ~new_G554_;
  assign new_G630_ = new_G540_ & new_G905_;
  assign new_G634_ = ~new_G540_ | ~new_G905_;
  assign new_G639_ = ~new_G636_;
  assign new_G642_ = ~new_G3082_ | ~new_G3085_;
  assign new_G3086_ = ~new_G3082_;
  assign new_G644_ = new_G460_ & new_G636_;
  assign new_G646_ = ~new_G3098_ | ~new_G3101_;
  assign new_G3102_ = ~new_G3098_;
  assign new_G654_ = ~G87 | ~new_G626_;
  assign new_G660_ = ~new_G657_;
  assign new_G678_ = ~new_G675_;
  assign new_G804_ = ~new_G860_ | ~new_G776_;
  assign new_G806_ = ~new_G860_ | ~new_G780_;
  assign new_G855_ = ~new_G736_ | ~new_G707_ | ~new_G721_;
  assign new_G867_ = ~new_G794_ | ~new_G736_ | ~new_G707_ | ~new_G724_;
  assign new_G903_ = ~new_G3090_ | ~new_G3093_;
  assign new_G3094_ = ~new_G3090_;
  assign new_G912_ = ~new_G3106_ | ~new_G3109_;
  assign new_G3110_ = ~new_G3106_;
  assign new_G915_ = ~new_G861_;
  assign new_G927_ = ~new_G893_;
  assign new_G941_ = ~new_G864_;
  assign new_G977_ = new_G828_ & new_G974_;
  assign new_G978_ = G150 & new_G975_;
  assign new_G984_ = new_G833_ & new_G981_;
  assign new_G985_ = G159 & new_G982_;
  assign new_G991_ = G77 & new_G988_;
  assign new_G992_ = G50 & new_G989_;
  assign new_G998_ = new_G839_ & new_G995_;
  assign new_G999_ = new_G828_ & new_G996_;
  assign new_G1005_ = new_G845_ & new_G1002_;
  assign new_G1006_ = new_G833_ & new_G1003_;
  assign new_G1012_ = G107 & new_G1009_;
  assign new_G1013_ = G77 & new_G1010_;
  assign new_G1019_ = G116 & new_G1016_;
  assign new_G1020_ = new_G839_ & new_G1017_;
  assign new_G1026_ = G283 & new_G1023_;
  assign new_G1027_ = new_G845_ & new_G1024_;
  assign new_G1060_ = G200 & new_G1054_;
  assign new_G1063_ = new_G1048_ & new_G1054_;
  assign new_G1066_ = new_G1049_ & new_G1057_;
  assign new_G1069_ = new_G1050_ & new_G1057_;
  assign new_G1527_ = ~new_G784_ | ~new_G794_;
  assign new_G1530_ = ~new_G776_ | ~new_G794_;
  assign new_G1542_ = ~new_G1541_ | ~new_G707_ | ~new_G721_;
  assign new_G1563_ = ~new_G784_ | ~new_G724_ | ~new_G732_;
  assign new_G1572_ = ~new_G724_ | ~new_G784_;
  assign new_G1581_ = ~new_G1512_;
  assign new_G1585_ = ~new_G1512_;
  assign new_G1589_ = ~new_G1512_;
  assign new_G1593_ = ~new_G1512_;
  assign new_G1597_ = ~new_G1512_;
  assign new_G1601_ = ~new_G1512_;
  assign new_G1605_ = ~new_G1512_;
  assign new_G1716_ = ~new_G1681_;
  assign new_G1718_ = new_G1681_ & new_G1699_;
  assign new_G1723_ = ~new_G1681_;
  assign new_G1725_ = new_G1681_ & new_G1699_;
  assign new_G1730_ = ~new_G1681_;
  assign new_G1732_ = new_G1681_ & new_G1699_;
  assign new_G1737_ = ~new_G1681_;
  assign new_G1739_ = new_G1681_ & new_G1699_;
  assign new_G1744_ = ~new_G1681_;
  assign new_G1746_ = new_G1681_ & new_G1699_;
  assign new_G1751_ = ~new_G1681_;
  assign new_G1753_ = new_G1681_ & new_G1699_;
  assign new_G1758_ = ~new_G1681_;
  assign new_G1760_ = new_G1681_ & new_G1699_;
  assign new_G1765_ = ~new_G1681_;
  assign new_G1767_ = new_G1681_ & new_G1699_;
  assign new_G1852_ = new_G1834_ & new_G1773_;
  assign new_G1856_ = ~G50 & ~new_G1773_;
  assign new_G1870_ = ~new_G807_;
  assign new_G1902_ = new_G1834_ & new_G1773_;
  assign new_G1906_ = ~G58 & ~new_G1773_;
  assign new_G1920_ = ~new_G807_;
  assign new_G1953_ = new_G1834_ & new_G1773_;
  assign new_G1957_ = ~G68 & ~new_G1773_;
  assign new_G1971_ = ~new_G807_;
  assign new_G2003_ = new_G1834_ & new_G1773_;
  assign new_G2007_ = ~G77 & ~new_G1773_;
  assign new_G2021_ = ~new_G807_;
  assign new_G2058_ = new_G1834_ & new_G1773_;
  assign new_G2062_ = ~G87 & ~new_G1773_;
  assign new_G2076_ = ~new_G823_;
  assign new_G2110_ = new_G1834_ & new_G1773_;
  assign new_G2114_ = ~G97 & ~new_G1773_;
  assign new_G2128_ = ~new_G816_;
  assign new_G2163_ = new_G1834_ & new_G1773_;
  assign new_G2167_ = ~G107 & ~new_G1773_;
  assign new_G2181_ = ~new_G816_;
  assign new_G2215_ = new_G1834_ & new_G1773_;
  assign new_G2219_ = ~G116 & ~new_G1773_;
  assign new_G2233_ = ~new_G816_;
  assign new_G2285_ = new_G2278_ & G213;
  assign new_G2288_ = ~new_G2278_ | ~G213;
  assign new_G2289_ = G343 & new_G2278_ & G213;
  assign new_G2293_ = ~G343 | ~new_G2278_ | ~G213;
  assign new_G2298_ = G343 & new_G2278_ & G213;
  assign new_G2302_ = ~G343 | ~new_G2278_ | ~G213;
  assign new_G2877_ = new_G2874_;
  assign new_G2983_ = ~new_G2955_ | ~new_G2956_;
  assign new_G2986_ = ~new_G2965_ | ~new_G2966_;
  assign new_G3014_ = ~new_G3010_;
  assign new_G3015_ = ~new_G3010_ | ~new_G3013_;
  assign new_G3023_ = ~new_G3017_;
  assign new_G3024_ = ~new_G3020_;
  assign new_G3033_ = ~new_G3027_;
  assign new_G3034_ = ~new_G3030_;
  assign new_G3043_ = ~new_G3037_;
  assign new_G3044_ = ~new_G3040_;
  assign G355 = ~new_G354_;
  assign new_G643_ = ~new_G3079_ | ~new_G3086_;
  assign new_G647_ = ~new_G3095_ | ~new_G3102_;
  assign new_G680_ = new_G650_ & new_G675_;
  assign new_G904_ = ~new_G3087_ | ~new_G3094_;
  assign new_G913_ = ~new_G3103_ | ~new_G3110_;
  assign new_G920_ = new_G588_ & new_G915_;
  assign new_G979_ = new_G978_ | new_G976_ | new_G977_;
  assign new_G993_ = new_G992_ | new_G990_ | new_G991_;
  assign new_G1000_ = new_G999_ | new_G997_ | new_G998_;
  assign new_G1007_ = new_G1006_ | new_G1004_ | new_G1005_;
  assign new_G1021_ = new_G1020_ | new_G1018_ | new_G1019_;
  assign new_G1028_ = new_G1027_ | new_G1025_ | new_G1026_;
  assign new_G1719_ = G77 & new_G1716_;
  assign new_G1721_ = G223 & new_G1718_;
  assign new_G1726_ = G87 & new_G1723_;
  assign new_G1728_ = G226 & new_G1725_;
  assign new_G1733_ = G97 & new_G1730_;
  assign new_G1735_ = G232 & new_G1732_;
  assign new_G1740_ = G107 & new_G1737_;
  assign new_G1742_ = G238 & new_G1739_;
  assign new_G1747_ = G116 & new_G1744_;
  assign new_G1749_ = G244 & new_G1746_;
  assign new_G1754_ = G283 & new_G1751_;
  assign new_G1756_ = G250 & new_G1753_;
  assign new_G1761_ = G294 & new_G1758_;
  assign new_G1763_ = G257 & new_G1760_;
  assign new_G1768_ = G303 & new_G1765_;
  assign new_G1770_ = G264 & new_G1767_;
  assign new_G1794_ = new_G1791_;
  assign new_G1799_ = ~new_G1791_;
  assign new_G1812_ = new_G1809_;
  assign new_G1817_ = ~new_G1809_;
  assign new_G1859_ = new_G1852_ & G50 & new_G1829_;
  assign new_G1909_ = new_G1902_ & G58 & new_G1829_;
  assign new_G1960_ = new_G1953_ & G68 & new_G1829_;
  assign new_G2010_ = new_G2003_ & G77 & new_G1829_;
  assign new_G2065_ = new_G2058_ & G87 & new_G2052_;
  assign new_G2117_ = new_G2110_ & G97 & new_G2052_;
  assign new_G2170_ = new_G2163_ & G107 & new_G2052_;
  assign new_G2222_ = new_G2215_ & G116 & new_G2052_;
  assign new_G2678_ = ~new_G956_;
  assign new_G2697_ = ~new_G956_;
  assign new_G2716_ = ~new_G956_;
  assign new_G2733_ = ~new_G956_;
  assign new_G2751_ = ~new_G956_;
  assign new_G2768_ = ~new_G956_;
  assign new_G2785_ = ~new_G956_;
  assign new_G2802_ = ~new_G956_;
  assign new_G3016_ = ~new_G3007_ | ~new_G3014_;
  assign new_G3025_ = ~new_G3020_ | ~new_G3023_;
  assign new_G3026_ = ~new_G3017_ | ~new_G3024_;
  assign new_G3035_ = ~new_G3030_ | ~new_G3033_;
  assign new_G3036_ = ~new_G3027_ | ~new_G3034_;
  assign new_G3045_ = ~new_G3040_ | ~new_G3043_;
  assign new_G3046_ = ~new_G3037_ | ~new_G3044_;
  assign new_G2989_ = ~new_G2983_;
  assign new_G2990_ = ~new_G2986_;
  assign new_G610_ = ~new_G804_;
  assign new_G613_ = new_G804_ & new_G806_;
  assign new_G616_ = ~new_G806_;
  assign new_G640_ = ~new_G642_ | ~new_G643_;
  assign new_G648_ = ~new_G646_ | ~new_G647_;
  assign new_G655_ = G58 & new_G442_ & new_G630_ & new_G635_;
  assign new_G665_ = ~new_G804_;
  assign new_G668_ = new_G804_ & new_G806_;
  assign new_G671_ = ~new_G806_;
  assign new_G683_ = ~new_G804_;
  assign new_G685_ = ~new_G806_;
  assign new_G688_ = new_G804_ & new_G806_;
  assign new_G694_ = ~new_G804_;
  assign new_G696_ = ~new_G806_;
  assign new_G699_ = new_G804_ & new_G806_;
  assign new_G870_ = new_G867_;
  assign new_G887_ = new_G867_;
  assign new_G901_ = ~new_G903_ | ~new_G904_;
  assign new_G910_ = ~new_G912_ | ~new_G913_;
  assign new_G914_ = ~new_G855_;
  assign new_G916_ = new_G855_ & new_G861_;
  assign new_G942_ = ~new_G855_;
  assign new_G943_ = new_G864_ & new_G855_;
  assign new_G1072_ = ~new_G1043_ | ~new_G1069_;
  assign new_G1084_ = ~new_G1043_ | ~new_G1066_;
  assign new_G1096_ = ~new_G1038_ | ~new_G1069_;
  assign new_G1108_ = ~new_G1038_ | ~new_G1066_;
  assign new_G1120_ = ~new_G1043_ | ~new_G1063_;
  assign new_G1132_ = ~new_G1043_ | ~new_G1060_;
  assign new_G1144_ = ~new_G1038_ | ~new_G1063_;
  assign new_G1156_ = ~new_G1038_ | ~new_G1060_;
  assign new_G1533_ = ~new_G1527_;
  assign new_G1534_ = ~new_G1530_;
  assign new_G1535_ = new_G1527_ & new_G1530_;
  assign new_G1545_ = new_G1542_;
  assign new_G1554_ = new_G1542_;
  assign new_G1610_ = ~new_G1572_;
  assign new_G1619_ = ~new_G1572_;
  assign new_G1628_ = ~new_G1572_;
  assign new_G1637_ = ~new_G1572_;
  assign new_G1646_ = ~new_G1563_;
  assign new_G1655_ = ~new_G1563_;
  assign new_G1664_ = ~new_G1563_;
  assign new_G1673_ = ~new_G1563_;
  assign new_G1722_ = new_G1721_ | new_G1719_ | new_G1720_;
  assign new_G1729_ = new_G1728_ | new_G1726_ | new_G1727_;
  assign new_G1736_ = new_G1735_ | new_G1733_ | new_G1734_;
  assign new_G1743_ = new_G1742_ | new_G1740_ | new_G1741_;
  assign new_G1750_ = new_G1749_ | new_G1747_ | new_G1748_;
  assign new_G1757_ = new_G1756_ | new_G1754_ | new_G1755_;
  assign new_G1764_ = new_G1763_ | new_G1761_ | new_G1762_;
  assign new_G1771_ = new_G1770_ | new_G1768_ | new_G1769_;
  assign new_G1853_ = new_G979_ & new_G1851_;
  assign new_G1954_ = new_G993_ & new_G1952_;
  assign new_G2004_ = new_G1000_ & new_G2002_;
  assign new_G2059_ = new_G1007_ & new_G2057_;
  assign new_G2164_ = new_G1021_ & new_G2162_;
  assign new_G2216_ = new_G1028_ & new_G2214_;
  assign new_G2485_ = new_G2293_;
  assign new_G2900_ = new_G2877_ & G2897;
  assign new_G2903_ = ~new_G2877_ | ~G2897;
  assign new_G2967_ = new_G557_;
  assign new_G2970_ = new_G562_;
  assign new_G2975_ = new_G557_;
  assign new_G2978_ = new_G562_;
  assign new_G3047_ = ~new_G3015_ | ~new_G3016_;
  assign new_G3050_ = ~new_G3025_ | ~new_G3026_;
  assign new_G3055_ = ~new_G3035_ | ~new_G3036_;
  assign new_G3058_ = ~new_G3045_ | ~new_G3046_;
  assign new_G574_ = ~new_G2986_ | ~new_G2989_;
  assign new_G575_ = ~new_G2983_ | ~new_G2990_;
  assign new_G617_ = new_G501_ & new_G613_;
  assign new_G641_ = new_G639_ & new_G640_ & new_G476_;
  assign new_G649_ = new_G530_ & new_G648_;
  assign new_G662_ = new_G655_ & new_G657_;
  assign new_G672_ = new_G513_ & new_G668_;
  assign new_G690_ = new_G654_ & new_G685_;
  assign new_G691_ = new_G540_ & new_G688_;
  assign new_G701_ = new_G634_ & new_G696_;
  assign new_G702_ = new_G526_ & new_G699_;
  assign new_G902_ = ~new_G901_;
  assign new_G911_ = ~new_G910_;
  assign new_G917_ = new_G650_ & new_G914_;
  assign new_G923_ = new_G586_ & new_G916_;
  assign new_G1538_ = new_G442_ & new_G1535_;
  assign new_G1871_ = new_G1870_ & new_G1817_ & G226;
  assign new_G1872_ = new_G807_ & new_G1817_ & G274;
  assign new_G1873_ = new_G1812_ & new_G1722_;
  assign new_G1921_ = new_G1920_ & new_G1817_ & G232;
  assign new_G1922_ = new_G807_ & new_G1817_ & G274;
  assign new_G1923_ = new_G1812_ & new_G1729_;
  assign new_G1972_ = new_G1971_ & new_G1817_ & G238;
  assign new_G1973_ = new_G807_ & new_G1817_ & G274;
  assign new_G1974_ = new_G1812_ & new_G1736_;
  assign new_G2022_ = new_G2021_ & new_G1817_ & G244;
  assign new_G2023_ = new_G807_ & new_G1817_ & G274;
  assign new_G2024_ = new_G1812_ & new_G1743_;
  assign new_G2077_ = new_G2076_ & new_G1799_ & G250;
  assign new_G2078_ = new_G823_ & new_G1799_ & G274;
  assign new_G2079_ = new_G1794_ & new_G1750_;
  assign new_G2129_ = new_G2128_ & new_G1799_ & G257;
  assign new_G2130_ = new_G816_ & new_G1799_ & G274;
  assign new_G2131_ = new_G1794_ & new_G1757_;
  assign new_G2182_ = new_G2181_ & new_G1799_ & G264;
  assign new_G2183_ = new_G816_ & new_G1799_ & G274;
  assign new_G2184_ = new_G1794_ & new_G1764_;
  assign new_G2234_ = new_G2233_ & new_G1799_ & G270;
  assign new_G2235_ = new_G816_ & new_G1799_ & G274;
  assign new_G2236_ = new_G1794_ & new_G1771_;
  assign new_G2973_ = ~new_G2967_;
  assign new_G2974_ = ~new_G2970_;
  assign new_G2981_ = ~new_G2975_;
  assign new_G2982_ = ~new_G2978_;
  assign new_G576_ = ~new_G574_ | ~new_G575_;
  assign new_G3053_ = ~new_G3047_;
  assign new_G3054_ = ~new_G3050_;
  assign new_G3061_ = ~new_G3055_;
  assign new_G3062_ = ~new_G3058_;
  assign new_G645_ = new_G641_ | new_G644_;
  assign new_G926_ = ~new_G887_;
  assign new_G928_ = new_G887_ & new_G893_;
  assign new_G947_ = new_G649_ & new_G942_;
  assign new_G983_ = new_G902_ & new_G980_;
  assign new_G1011_ = new_G911_ & new_G1008_;
  assign new_G1075_ = new_G1072_;
  assign new_G1087_ = new_G1084_;
  assign new_G1099_ = new_G1096_;
  assign new_G1111_ = new_G1108_;
  assign new_G1123_ = new_G1120_;
  assign new_G1135_ = new_G1132_;
  assign new_G1147_ = new_G1144_;
  assign new_G1159_ = new_G1156_;
  assign new_G1168_ = new_G1072_;
  assign new_G1177_ = new_G1084_;
  assign new_G1186_ = new_G1096_;
  assign new_G1195_ = new_G1108_;
  assign new_G1204_ = new_G1120_;
  assign new_G1213_ = new_G1132_;
  assign new_G1222_ = new_G1144_;
  assign new_G1231_ = new_G1156_;
  assign new_G1609_ = ~new_G1545_;
  assign new_G1611_ = new_G1545_ & new_G1572_;
  assign new_G1618_ = ~new_G1545_;
  assign new_G1620_ = new_G1545_ & new_G1572_;
  assign new_G1627_ = ~new_G1545_;
  assign new_G1629_ = new_G1545_ & new_G1572_;
  assign new_G1636_ = ~new_G1545_;
  assign new_G1638_ = new_G1545_ & new_G1572_;
  assign new_G1645_ = ~new_G1554_;
  assign new_G1647_ = new_G1554_ & new_G1563_;
  assign new_G1654_ = ~new_G1554_;
  assign new_G1656_ = new_G1554_ & new_G1563_;
  assign new_G1663_ = ~new_G1554_;
  assign new_G1665_ = new_G1554_ & new_G1563_;
  assign new_G1672_ = ~new_G1554_;
  assign new_G1674_ = new_G1554_ & new_G1563_;
  assign new_G1862_ = new_G1859_ | new_G1853_ | new_G1856_;
  assign new_G1866_ = ~new_G1859_ & ~new_G1853_ & ~new_G1856_;
  assign new_G1874_ = new_G1873_ | new_G1871_ | new_G1872_;
  assign new_G1924_ = new_G1923_ | new_G1921_ | new_G1922_;
  assign new_G1963_ = new_G1960_ | new_G1954_ | new_G1957_;
  assign new_G1967_ = ~new_G1960_ & ~new_G1954_ & ~new_G1957_;
  assign new_G1975_ = new_G1974_ | new_G1972_ | new_G1973_;
  assign new_G2013_ = new_G2010_ | new_G2004_ | new_G2007_;
  assign new_G2017_ = ~new_G2010_ & ~new_G2004_ & ~new_G2007_;
  assign new_G2025_ = new_G2024_ | new_G2022_ | new_G2023_;
  assign new_G2068_ = new_G2065_ | new_G2059_ | new_G2062_;
  assign new_G2072_ = ~new_G2065_ & ~new_G2059_ & ~new_G2062_;
  assign new_G2080_ = new_G2079_ | new_G2077_ | new_G2078_;
  assign new_G2132_ = new_G2131_ | new_G2129_ | new_G2130_;
  assign new_G2173_ = new_G2170_ | new_G2164_ | new_G2167_;
  assign new_G2177_ = ~new_G2170_ & ~new_G2164_ & ~new_G2167_;
  assign new_G2185_ = new_G2184_ | new_G2182_ | new_G2183_;
  assign new_G2225_ = new_G2222_ | new_G2216_ | new_G2219_;
  assign new_G2229_ = ~new_G2222_ & ~new_G2216_ & ~new_G2219_;
  assign new_G2237_ = new_G2236_ | new_G2234_ | new_G2235_;
  assign new_G2488_ = ~new_G2485_;
  assign new_G2679_ = ~new_G870_;
  assign new_G2680_ = new_G956_ & new_G870_;
  assign new_G2698_ = ~new_G870_;
  assign new_G2699_ = new_G956_ & new_G870_;
  assign new_G2717_ = ~new_G870_;
  assign new_G2718_ = new_G956_ & new_G870_;
  assign new_G2734_ = ~new_G870_;
  assign new_G2735_ = new_G956_ & new_G870_;
  assign new_G2752_ = ~new_G870_;
  assign new_G2753_ = new_G956_ & new_G870_;
  assign new_G2769_ = ~new_G870_;
  assign new_G2770_ = new_G956_ & new_G870_;
  assign new_G2786_ = ~new_G870_;
  assign new_G2787_ = new_G956_ & new_G870_;
  assign new_G2803_ = ~new_G870_;
  assign new_G2804_ = new_G956_ & new_G870_;
  assign new_G359_ = new_G923_ | new_G917_ | new_G920_;
  assign new_G1029_ = ~new_G923_ & ~new_G917_ & ~new_G920_;
  assign new_G565_ = ~new_G2970_ | ~new_G2973_;
  assign new_G566_ = ~new_G2967_ | ~new_G2974_;
  assign new_G569_ = ~new_G2978_ | ~new_G2981_;
  assign new_G570_ = ~new_G2975_ | ~new_G2982_;
  assign new_G589_ = ~new_G3050_ | ~new_G3053_;
  assign new_G590_ = ~new_G3047_ | ~new_G3054_;
  assign new_G595_ = ~new_G3058_ | ~new_G3061_;
  assign new_G596_ = ~new_G3055_ | ~new_G3062_;
  assign new_G929_ = new_G650_ & new_G926_;
  assign new_G938_ = new_G630_ & new_G928_;
  assign new_G944_ = new_G645_ & new_G941_;
  assign new_G986_ = new_G985_ | new_G983_ | new_G984_;
  assign new_G1014_ = new_G1013_ | new_G1011_ | new_G1012_;
  assign new_G1616_ = new_G442_ & new_G1611_;
  assign new_G1625_ = new_G456_ & new_G1620_;
  assign new_G1634_ = new_G463_ & new_G1629_;
  assign new_G1643_ = new_G479_ & new_G1638_;
  assign new_G360_ = ~new_G1029_;
  assign new_G567_ = ~new_G565_ | ~new_G566_;
  assign new_G571_ = ~new_G569_ | ~new_G570_;
  assign new_G579_ = new_G576_;
  assign new_G591_ = ~new_G589_ | ~new_G590_;
  assign new_G597_ = ~new_G595_ | ~new_G596_;
  assign new_G614_ = new_G576_ & new_G610_;
  assign new_G1240_ = ~new_G1075_;
  assign new_G1241_ = ~new_G1087_;
  assign new_G1242_ = ~new_G1099_;
  assign new_G1243_ = ~new_G1111_;
  assign new_G1244_ = ~new_G1123_;
  assign new_G1245_ = ~new_G1135_;
  assign new_G1246_ = ~new_G1147_;
  assign new_G1247_ = ~new_G1159_;
  assign new_G1257_ = ~new_G1075_;
  assign new_G1258_ = ~new_G1087_;
  assign new_G1259_ = ~new_G1099_;
  assign new_G1260_ = ~new_G1111_;
  assign new_G1261_ = ~new_G1123_;
  assign new_G1262_ = ~new_G1135_;
  assign new_G1263_ = ~new_G1147_;
  assign new_G1264_ = ~new_G1159_;
  assign new_G1274_ = ~new_G1075_;
  assign new_G1275_ = ~new_G1087_;
  assign new_G1276_ = ~new_G1099_;
  assign new_G1277_ = ~new_G1111_;
  assign new_G1278_ = ~new_G1123_;
  assign new_G1279_ = ~new_G1135_;
  assign new_G1280_ = ~new_G1147_;
  assign new_G1281_ = ~new_G1159_;
  assign new_G1291_ = ~new_G1075_;
  assign new_G1292_ = ~new_G1087_;
  assign new_G1293_ = ~new_G1099_;
  assign new_G1294_ = ~new_G1111_;
  assign new_G1295_ = ~new_G1123_;
  assign new_G1296_ = ~new_G1135_;
  assign new_G1297_ = ~new_G1147_;
  assign new_G1298_ = ~new_G1159_;
  assign new_G1308_ = ~new_G1075_;
  assign new_G1309_ = ~new_G1087_;
  assign new_G1310_ = ~new_G1099_;
  assign new_G1311_ = ~new_G1111_;
  assign new_G1312_ = ~new_G1123_;
  assign new_G1313_ = ~new_G1135_;
  assign new_G1314_ = ~new_G1147_;
  assign new_G1315_ = ~new_G1159_;
  assign new_G1325_ = ~new_G1075_;
  assign new_G1326_ = ~new_G1087_;
  assign new_G1327_ = ~new_G1099_;
  assign new_G1328_ = ~new_G1111_;
  assign new_G1329_ = ~new_G1123_;
  assign new_G1330_ = ~new_G1135_;
  assign new_G1331_ = ~new_G1147_;
  assign new_G1332_ = ~new_G1159_;
  assign new_G1342_ = ~new_G1075_;
  assign new_G1343_ = ~new_G1087_;
  assign new_G1344_ = ~new_G1099_;
  assign new_G1345_ = ~new_G1111_;
  assign new_G1346_ = ~new_G1123_;
  assign new_G1347_ = ~new_G1135_;
  assign new_G1348_ = ~new_G1147_;
  assign new_G1349_ = ~new_G1159_;
  assign new_G1359_ = ~new_G1075_;
  assign new_G1360_ = ~new_G1087_;
  assign new_G1361_ = ~new_G1099_;
  assign new_G1362_ = ~new_G1111_;
  assign new_G1363_ = ~new_G1123_;
  assign new_G1364_ = ~new_G1135_;
  assign new_G1365_ = ~new_G1147_;
  assign new_G1366_ = ~new_G1159_;
  assign new_G1376_ = ~new_G1168_;
  assign new_G1377_ = ~new_G1177_;
  assign new_G1378_ = ~new_G1186_;
  assign new_G1379_ = ~new_G1195_;
  assign new_G1380_ = ~new_G1204_;
  assign new_G1381_ = ~new_G1213_;
  assign new_G1382_ = ~new_G1222_;
  assign new_G1383_ = ~new_G1231_;
  assign new_G1393_ = ~new_G1168_;
  assign new_G1394_ = ~new_G1177_;
  assign new_G1395_ = ~new_G1186_;
  assign new_G1396_ = ~new_G1195_;
  assign new_G1397_ = ~new_G1204_;
  assign new_G1398_ = ~new_G1213_;
  assign new_G1399_ = ~new_G1222_;
  assign new_G1400_ = ~new_G1231_;
  assign new_G1410_ = ~new_G1168_;
  assign new_G1411_ = ~new_G1177_;
  assign new_G1412_ = ~new_G1186_;
  assign new_G1413_ = ~new_G1195_;
  assign new_G1414_ = ~new_G1204_;
  assign new_G1415_ = ~new_G1213_;
  assign new_G1416_ = ~new_G1222_;
  assign new_G1417_ = ~new_G1231_;
  assign new_G1427_ = ~new_G1168_;
  assign new_G1428_ = ~new_G1177_;
  assign new_G1429_ = ~new_G1186_;
  assign new_G1430_ = ~new_G1195_;
  assign new_G1431_ = ~new_G1204_;
  assign new_G1432_ = ~new_G1213_;
  assign new_G1433_ = ~new_G1222_;
  assign new_G1434_ = ~new_G1231_;
  assign new_G1444_ = ~new_G1168_;
  assign new_G1445_ = ~new_G1177_;
  assign new_G1446_ = ~new_G1186_;
  assign new_G1447_ = ~new_G1195_;
  assign new_G1448_ = ~new_G1204_;
  assign new_G1449_ = ~new_G1213_;
  assign new_G1450_ = ~new_G1222_;
  assign new_G1451_ = ~new_G1231_;
  assign new_G1461_ = ~new_G1168_;
  assign new_G1462_ = ~new_G1177_;
  assign new_G1463_ = ~new_G1186_;
  assign new_G1464_ = ~new_G1195_;
  assign new_G1465_ = ~new_G1204_;
  assign new_G1466_ = ~new_G1213_;
  assign new_G1467_ = ~new_G1222_;
  assign new_G1468_ = ~new_G1231_;
  assign new_G1478_ = ~new_G1168_;
  assign new_G1479_ = ~new_G1177_;
  assign new_G1480_ = ~new_G1186_;
  assign new_G1481_ = ~new_G1195_;
  assign new_G1482_ = ~new_G1204_;
  assign new_G1483_ = ~new_G1213_;
  assign new_G1484_ = ~new_G1222_;
  assign new_G1485_ = ~new_G1231_;
  assign new_G1495_ = ~new_G1168_;
  assign new_G1496_ = ~new_G1177_;
  assign new_G1497_ = ~new_G1186_;
  assign new_G1498_ = ~new_G1195_;
  assign new_G1499_ = ~new_G1204_;
  assign new_G1500_ = ~new_G1213_;
  assign new_G1501_ = ~new_G1222_;
  assign new_G1502_ = ~new_G1231_;
  assign new_G1877_ = new_G1874_;
  assign new_G1880_ = ~new_G1874_;
  assign new_G1891_ = ~new_G1866_;
  assign new_G1903_ = new_G986_ & new_G1901_;
  assign new_G1927_ = new_G1924_;
  assign new_G1930_ = ~new_G1924_;
  assign new_G1978_ = new_G1975_;
  assign new_G1981_ = ~new_G1975_;
  assign new_G1992_ = ~new_G1967_;
  assign new_G2028_ = new_G2025_;
  assign new_G2031_ = ~new_G2025_;
  assign new_G2042_ = ~new_G2017_;
  assign new_G2085_ = new_G2080_;
  assign new_G2088_ = ~new_G2080_;
  assign new_G2099_ = ~new_G2072_;
  assign new_G2111_ = new_G1014_ & new_G2109_;
  assign new_G2137_ = new_G2132_;
  assign new_G2140_ = ~new_G2132_;
  assign new_G2190_ = new_G2185_;
  assign new_G2193_ = ~new_G2185_;
  assign new_G2204_ = ~new_G2177_;
  assign new_G2242_ = new_G2237_;
  assign new_G2245_ = ~new_G2237_;
  assign new_G2256_ = ~new_G2229_;
  assign new_G2320_ = new_G2285_ & new_G1862_;
  assign new_G2341_ = new_G2289_ & new_G1963_;
  assign new_G2354_ = new_G2289_ & new_G2013_;
  assign new_G2367_ = new_G2289_ & new_G2068_;
  assign new_G2383_ = new_G2298_ & new_G2173_;
  assign new_G2391_ = new_G2298_ & new_G2225_;
  assign new_G2474_ = ~new_G2080_;
  assign new_G2475_ = ~new_G2132_;
  assign new_G2476_ = ~new_G2185_;
  assign new_G2477_ = ~new_G2237_;
  assign new_G2482_ = new_G2481_ & new_G2237_ & new_G2185_ & new_G2080_ & new_G2132_;
  assign G361 = ~new_G359_ | ~new_G360_;
  assign new_G568_ = ~new_G567_;
  assign new_G618_ = new_G617_ | new_G614_ | new_G616_;
  assign new_G1248_ = G124 & new_G1240_;
  assign new_G1249_ = G159 & new_G1241_;
  assign new_G1250_ = G150 & new_G1242_;
  assign new_G1251_ = G143 & new_G1243_;
  assign new_G1252_ = G137 & new_G1244_;
  assign new_G1253_ = G132 & new_G1245_;
  assign new_G1254_ = G128 & new_G1246_;
  assign new_G1255_ = G125 & new_G1247_;
  assign new_G1265_ = G125 & new_G1257_;
  assign new_G1266_ = new_G432_ & new_G1258_;
  assign new_G1267_ = G159 & new_G1259_;
  assign new_G1268_ = G150 & new_G1260_;
  assign new_G1269_ = G143 & new_G1261_;
  assign new_G1270_ = G137 & new_G1262_;
  assign new_G1271_ = G132 & new_G1263_;
  assign new_G1272_ = G128 & new_G1264_;
  assign new_G1282_ = G128 & new_G1274_;
  assign new_G1283_ = new_G447_ & new_G1275_;
  assign new_G1284_ = new_G432_ & new_G1276_;
  assign new_G1285_ = G159 & new_G1277_;
  assign new_G1286_ = G150 & new_G1278_;
  assign new_G1287_ = G143 & new_G1279_;
  assign new_G1288_ = G137 & new_G1280_;
  assign new_G1289_ = G132 & new_G1281_;
  assign new_G1299_ = G132 & new_G1291_;
  assign new_G1300_ = new_G467_ & new_G1292_;
  assign new_G1301_ = new_G447_ & new_G1293_;
  assign new_G1302_ = new_G432_ & new_G1294_;
  assign new_G1303_ = G159 & new_G1295_;
  assign new_G1304_ = G150 & new_G1296_;
  assign new_G1305_ = G143 & new_G1297_;
  assign new_G1306_ = G137 & new_G1298_;
  assign new_G1316_ = G137 & new_G1308_;
  assign new_G1317_ = new_G483_ & new_G1309_;
  assign new_G1318_ = new_G467_ & new_G1310_;
  assign new_G1319_ = new_G447_ & new_G1311_;
  assign new_G1320_ = new_G432_ & new_G1312_;
  assign new_G1321_ = G159 & new_G1313_;
  assign new_G1322_ = G150 & new_G1314_;
  assign new_G1323_ = G143 & new_G1315_;
  assign new_G1333_ = G143 & new_G1325_;
  assign new_G1334_ = new_G492_ & new_G1326_;
  assign new_G1335_ = new_G483_ & new_G1327_;
  assign new_G1336_ = new_G467_ & new_G1328_;
  assign new_G1337_ = new_G447_ & new_G1329_;
  assign new_G1338_ = new_G432_ & new_G1330_;
  assign new_G1339_ = G159 & new_G1331_;
  assign new_G1340_ = G150 & new_G1332_;
  assign new_G1350_ = G150 & new_G1342_;
  assign new_G1351_ = new_G504_ & new_G1343_;
  assign new_G1352_ = new_G492_ & new_G1344_;
  assign new_G1353_ = new_G483_ & new_G1345_;
  assign new_G1354_ = new_G467_ & new_G1346_;
  assign new_G1355_ = new_G447_ & new_G1347_;
  assign new_G1356_ = new_G432_ & new_G1348_;
  assign new_G1357_ = G159 & new_G1349_;
  assign new_G1367_ = G159 & new_G1359_;
  assign new_G1368_ = new_G517_ & new_G1360_;
  assign new_G1369_ = new_G504_ & new_G1361_;
  assign new_G1370_ = new_G492_ & new_G1362_;
  assign new_G1371_ = new_G483_ & new_G1363_;
  assign new_G1372_ = new_G467_ & new_G1364_;
  assign new_G1373_ = new_G447_ & new_G1365_;
  assign new_G1374_ = new_G432_ & new_G1366_;
  assign new_G1384_ = G283 & new_G1376_;
  assign new_G1385_ = new_G447_ & new_G1377_;
  assign new_G1386_ = new_G467_ & new_G1378_;
  assign new_G1387_ = new_G483_ & new_G1379_;
  assign new_G1388_ = new_G492_ & new_G1380_;
  assign new_G1389_ = new_G504_ & new_G1381_;
  assign new_G1390_ = new_G517_ & new_G1382_;
  assign new_G1391_ = new_G530_ & new_G1383_;
  assign new_G1401_ = G294 & new_G1393_;
  assign new_G1402_ = new_G467_ & new_G1394_;
  assign new_G1403_ = new_G483_ & new_G1395_;
  assign new_G1404_ = new_G492_ & new_G1396_;
  assign new_G1405_ = new_G504_ & new_G1397_;
  assign new_G1406_ = new_G517_ & new_G1398_;
  assign new_G1407_ = new_G530_ & new_G1399_;
  assign new_G1408_ = G283 & new_G1400_;
  assign new_G1418_ = G303 & new_G1410_;
  assign new_G1419_ = new_G483_ & new_G1411_;
  assign new_G1420_ = new_G492_ & new_G1412_;
  assign new_G1421_ = new_G504_ & new_G1413_;
  assign new_G1422_ = new_G517_ & new_G1414_;
  assign new_G1423_ = new_G530_ & new_G1415_;
  assign new_G1424_ = G283 & new_G1416_;
  assign new_G1425_ = G294 & new_G1417_;
  assign new_G1435_ = G311 & new_G1427_;
  assign new_G1436_ = new_G492_ & new_G1428_;
  assign new_G1437_ = new_G504_ & new_G1429_;
  assign new_G1438_ = new_G517_ & new_G1430_;
  assign new_G1439_ = new_G530_ & new_G1431_;
  assign new_G1440_ = G283 & new_G1432_;
  assign new_G1441_ = G294 & new_G1433_;
  assign new_G1442_ = G303 & new_G1434_;
  assign new_G1452_ = G317 & new_G1444_;
  assign new_G1453_ = new_G504_ & new_G1445_;
  assign new_G1454_ = new_G517_ & new_G1446_;
  assign new_G1455_ = new_G530_ & new_G1447_;
  assign new_G1456_ = G283 & new_G1448_;
  assign new_G1457_ = G294 & new_G1449_;
  assign new_G1458_ = G303 & new_G1450_;
  assign new_G1459_ = G311 & new_G1451_;
  assign new_G1469_ = G322 & new_G1461_;
  assign new_G1470_ = new_G517_ & new_G1462_;
  assign new_G1471_ = new_G530_ & new_G1463_;
  assign new_G1472_ = G283 & new_G1464_;
  assign new_G1473_ = G294 & new_G1465_;
  assign new_G1474_ = G303 & new_G1466_;
  assign new_G1475_ = G311 & new_G1467_;
  assign new_G1476_ = G317 & new_G1468_;
  assign new_G1486_ = G326 & new_G1478_;
  assign new_G1487_ = new_G530_ & new_G1479_;
  assign new_G1488_ = G283 & new_G1480_;
  assign new_G1489_ = G294 & new_G1481_;
  assign new_G1490_ = G303 & new_G1482_;
  assign new_G1491_ = G311 & new_G1483_;
  assign new_G1492_ = G317 & new_G1484_;
  assign new_G1493_ = G322 & new_G1485_;
  assign new_G1503_ = G329 & new_G1495_;
  assign new_G1504_ = G283 & new_G1496_;
  assign new_G1505_ = G294 & new_G1497_;
  assign new_G1506_ = G303 & new_G1498_;
  assign new_G1507_ = G311 & new_G1499_;
  assign new_G1508_ = G317 & new_G1500_;
  assign new_G1509_ = G322 & new_G1501_;
  assign new_G1510_ = G326 & new_G1502_;
  assign new_G2483_ = new_G2478_ & new_G2477_ & new_G2476_ & new_G2474_ & new_G2475_;
  assign new_G600_ = new_G597_;
  assign new_G661_ = new_G568_ & new_G660_;
  assign new_G669_ = new_G597_ & new_G665_;
  assign new_G679_ = new_G591_ & new_G678_;
  assign new_G1256_ = ~new_G1255_ & ~new_G1254_ & ~new_G1253_ & ~new_G1252_ & ~new_G1251_ & ~new_G1250_ & ~new_G1248_ & ~new_G1249_;
  assign new_G1273_ = ~new_G1272_ & ~new_G1271_ & ~new_G1270_ & ~new_G1269_ & ~new_G1268_ & ~new_G1267_ & ~new_G1265_ & ~new_G1266_;
  assign new_G1290_ = ~new_G1289_ & ~new_G1288_ & ~new_G1287_ & ~new_G1286_ & ~new_G1285_ & ~new_G1284_ & ~new_G1282_ & ~new_G1283_;
  assign new_G1307_ = ~new_G1306_ & ~new_G1305_ & ~new_G1304_ & ~new_G1303_ & ~new_G1302_ & ~new_G1301_ & ~new_G1299_ & ~new_G1300_;
  assign new_G1324_ = ~new_G1323_ & ~new_G1322_ & ~new_G1321_ & ~new_G1320_ & ~new_G1319_ & ~new_G1318_ & ~new_G1316_ & ~new_G1317_;
  assign new_G1341_ = ~new_G1340_ & ~new_G1339_ & ~new_G1338_ & ~new_G1337_ & ~new_G1336_ & ~new_G1335_ & ~new_G1333_ & ~new_G1334_;
  assign new_G1358_ = ~new_G1357_ & ~new_G1356_ & ~new_G1355_ & ~new_G1354_ & ~new_G1353_ & ~new_G1352_ & ~new_G1350_ & ~new_G1351_;
  assign new_G1375_ = ~new_G1374_ & ~new_G1373_ & ~new_G1372_ & ~new_G1371_ & ~new_G1370_ & ~new_G1369_ & ~new_G1367_ & ~new_G1368_;
  assign new_G1392_ = ~new_G1391_ & ~new_G1390_ & ~new_G1389_ & ~new_G1388_ & ~new_G1387_ & ~new_G1386_ & ~new_G1384_ & ~new_G1385_;
  assign new_G1409_ = ~new_G1408_ & ~new_G1407_ & ~new_G1406_ & ~new_G1405_ & ~new_G1404_ & ~new_G1403_ & ~new_G1401_ & ~new_G1402_;
  assign new_G1426_ = ~new_G1425_ & ~new_G1424_ & ~new_G1423_ & ~new_G1422_ & ~new_G1421_ & ~new_G1420_ & ~new_G1418_ & ~new_G1419_;
  assign new_G1443_ = ~new_G1442_ & ~new_G1441_ & ~new_G1440_ & ~new_G1439_ & ~new_G1438_ & ~new_G1437_ & ~new_G1435_ & ~new_G1436_;
  assign new_G1460_ = ~new_G1459_ & ~new_G1458_ & ~new_G1457_ & ~new_G1456_ & ~new_G1455_ & ~new_G1454_ & ~new_G1452_ & ~new_G1453_;
  assign new_G1477_ = ~new_G1476_ & ~new_G1475_ & ~new_G1474_ & ~new_G1473_ & ~new_G1472_ & ~new_G1471_ & ~new_G1469_ & ~new_G1470_;
  assign new_G1494_ = ~new_G1493_ & ~new_G1492_ & ~new_G1491_ & ~new_G1490_ & ~new_G1489_ & ~new_G1488_ & ~new_G1486_ & ~new_G1487_;
  assign new_G1511_ = ~new_G1510_ & ~new_G1509_ & ~new_G1508_ & ~new_G1507_ & ~new_G1506_ & ~new_G1505_ & ~new_G1503_ & ~new_G1504_;
  assign new_G1652_ = new_G618_ & new_G1647_;
  assign new_G1883_ = new_G1877_ & G169 & new_G1862_;
  assign new_G1886_ = new_G1880_ & G179 & new_G1862_;
  assign new_G1889_ = new_G1880_ & G190 & new_G1866_;
  assign new_G1890_ = new_G1877_ & G200 & new_G1866_;
  assign new_G1912_ = new_G1909_ | new_G1903_ | new_G1906_;
  assign new_G1916_ = ~new_G1909_ & ~new_G1903_ & ~new_G1906_;
  assign new_G1984_ = new_G1978_ & G169 & new_G1963_;
  assign new_G1987_ = new_G1981_ & G179 & new_G1963_;
  assign new_G1990_ = new_G1981_ & G190 & new_G1967_;
  assign new_G1991_ = new_G1978_ & G200 & new_G1967_;
  assign new_G2034_ = new_G2028_ & G169 & new_G2013_;
  assign new_G2037_ = new_G2031_ & G179 & new_G2013_;
  assign new_G2040_ = new_G2031_ & G190 & new_G2017_;
  assign new_G2041_ = new_G2028_ & G200 & new_G2017_;
  assign new_G2091_ = new_G2085_ & G169 & new_G2068_;
  assign new_G2094_ = new_G2088_ & G179 & new_G2068_;
  assign new_G2097_ = new_G2088_ & G190 & new_G2072_;
  assign new_G2098_ = new_G2085_ & G200 & new_G2072_;
  assign new_G2120_ = new_G2117_ | new_G2111_ | new_G2114_;
  assign new_G2124_ = ~new_G2117_ & ~new_G2111_ & ~new_G2114_;
  assign new_G2196_ = new_G2190_ & G169 & new_G2173_;
  assign new_G2199_ = new_G2193_ & G179 & new_G2173_;
  assign new_G2202_ = new_G2193_ & G190 & new_G2177_;
  assign new_G2203_ = new_G2190_ & G200 & new_G2177_;
  assign new_G2248_ = new_G2242_ & G169 & new_G2225_;
  assign new_G2251_ = new_G2245_ & G179 & new_G2225_;
  assign new_G2254_ = new_G2245_ & G190 & new_G2229_;
  assign new_G2255_ = new_G2242_ & G200 & new_G2229_;
  assign new_G2484_ = new_G2482_ | new_G2483_;
  assign new_G2991_ = new_G571_;
  assign new_G2994_ = new_G579_;
  assign new_G2999_ = new_G571_;
  assign new_G3002_ = new_G579_;
  assign new_G3063_ = new_G591_;
  assign new_G3071_ = new_G591_;
  assign new_G3124_ = new_G2320_;
  assign new_G3134_ = new_G2320_;
  assign new_G3158_ = new_G2341_;
  assign new_G3166_ = new_G2341_;
  assign new_G3174_ = new_G2354_;
  assign new_G3182_ = new_G2354_;
  assign new_G3190_ = new_G2367_;
  assign new_G3200_ = new_G2367_;
  assign new_G3224_ = new_G2383_;
  assign new_G3232_ = new_G2383_;
  assign new_G3240_ = new_G2391_;
  assign new_G3248_ = new_G2391_;
  assign new_G663_ = ~new_G661_ & ~new_G662_;
  assign new_G673_ = new_G672_ | new_G669_ | new_G671_;
  assign new_G681_ = ~new_G679_ & ~new_G680_;
  assign new_G1536_ = new_G1256_ & new_G1533_;
  assign new_G1537_ = new_G1392_ & new_G1534_;
  assign new_G1582_ = new_G1273_ & new_G1581_;
  assign new_G1583_ = new_G1409_ & new_G1512_;
  assign new_G1586_ = new_G1290_ & new_G1585_;
  assign new_G1587_ = new_G1426_ & new_G1512_;
  assign new_G1590_ = new_G1307_ & new_G1589_;
  assign new_G1591_ = new_G1443_ & new_G1512_;
  assign new_G1594_ = new_G1324_ & new_G1593_;
  assign new_G1595_ = new_G1460_ & new_G1512_;
  assign new_G1598_ = new_G1341_ & new_G1597_;
  assign new_G1599_ = new_G1477_ & new_G1512_;
  assign new_G1602_ = new_G1358_ & new_G1601_;
  assign new_G1603_ = new_G1494_ & new_G1512_;
  assign new_G1606_ = new_G1375_ & new_G1605_;
  assign new_G1607_ = new_G1511_ & new_G1512_;
  assign new_G1894_ = new_G1891_ | new_G1889_ | new_G1890_;
  assign new_G1997_ = new_G1992_ | new_G1990_ | new_G1991_;
  assign new_G2047_ = new_G2042_ | new_G2040_ | new_G2041_;
  assign new_G2102_ = new_G2099_ | new_G2097_ | new_G2098_;
  assign new_G2209_ = new_G2204_ | new_G2202_ | new_G2203_;
  assign new_G2261_ = new_G2256_ | new_G2254_ | new_G2255_;
  assign new_G2489_ = new_G2484_ & new_G2488_;
  assign new_G3005_ = ~new_G2999_;
  assign new_G3006_ = ~new_G3002_;
  assign new_G3077_ = ~new_G3071_;
  assign new_G3069_ = ~new_G3063_;
  assign new_G2997_ = ~new_G2991_;
  assign new_G2998_ = ~new_G2994_;
  assign new_G689_ = new_G681_ & new_G683_;
  assign new_G700_ = new_G663_ & new_G694_;
  assign new_G1539_ = new_G1538_ | new_G1536_ | new_G1537_;
  assign new_G1584_ = new_G1582_ | new_G1583_;
  assign new_G1588_ = new_G1586_ | new_G1587_;
  assign new_G1592_ = new_G1590_ | new_G1591_;
  assign new_G1596_ = new_G1594_ | new_G1595_;
  assign new_G1600_ = new_G1598_ | new_G1599_;
  assign new_G1604_ = new_G1602_ | new_G1603_;
  assign new_G1608_ = new_G1606_ | new_G1607_;
  assign new_G1661_ = new_G673_ & new_G1656_;
  assign new_G1892_ = new_G1883_ | new_G1886_;
  assign new_G1893_ = ~new_G1883_ & ~new_G1886_;
  assign new_G1933_ = new_G1927_ & G169 & new_G1912_;
  assign new_G1936_ = new_G1930_ & G179 & new_G1912_;
  assign new_G1939_ = new_G1930_ & G190 & new_G1916_;
  assign new_G1940_ = new_G1927_ & G200 & new_G1916_;
  assign new_G1941_ = ~new_G1916_;
  assign new_G1993_ = new_G1984_ | new_G1987_;
  assign new_G1996_ = ~new_G1984_ & ~new_G1987_;
  assign new_G2043_ = new_G2034_ | new_G2037_;
  assign new_G2046_ = ~new_G2034_ & ~new_G2037_;
  assign new_G2100_ = new_G2091_ | new_G2094_;
  assign new_G2101_ = ~new_G2091_ & ~new_G2094_;
  assign new_G2143_ = new_G2137_ & G169 & new_G2120_;
  assign new_G2146_ = new_G2140_ & G179 & new_G2120_;
  assign new_G2149_ = new_G2140_ & G190 & new_G2124_;
  assign new_G2150_ = new_G2137_ & G200 & new_G2124_;
  assign new_G2151_ = ~new_G2124_;
  assign new_G2205_ = new_G2196_ | new_G2199_;
  assign new_G2208_ = ~new_G2196_ & ~new_G2199_;
  assign new_G2257_ = new_G2248_ | new_G2251_;
  assign new_G2260_ = ~new_G2248_ & ~new_G2251_;
  assign new_G3138_ = ~new_G3134_;
  assign new_G2328_ = new_G2285_ & new_G1912_;
  assign new_G3162_ = ~new_G3158_;
  assign new_G3170_ = ~new_G3166_;
  assign new_G3178_ = ~new_G3174_;
  assign new_G3186_ = ~new_G3182_;
  assign new_G3204_ = ~new_G3200_;
  assign new_G2375_ = new_G2298_ & new_G2120_;
  assign new_G3236_ = ~new_G3232_;
  assign new_G3244_ = ~new_G3240_;
  assign new_G3252_ = ~new_G3248_;
  assign new_G3228_ = ~new_G3224_;
  assign new_G3066_ = new_G600_;
  assign new_G3074_ = new_G600_;
  assign new_G3128_ = ~new_G3124_;
  assign new_G3194_ = ~new_G3190_;
  assign new_G619_ = ~new_G2994_ | ~new_G2997_;
  assign new_G620_ = ~new_G2991_ | ~new_G2998_;
  assign new_G582_ = ~new_G3002_ | ~new_G3005_;
  assign new_G583_ = ~new_G2999_ | ~new_G3006_;
  assign new_G692_ = new_G691_ | new_G689_ | new_G690_;
  assign new_G703_ = new_G702_ | new_G700_ | new_G701_;
  assign new_G1612_ = new_G1539_ & new_G1609_;
  assign new_G1621_ = new_G1584_ & new_G1618_;
  assign new_G1630_ = new_G1588_ & new_G1627_;
  assign new_G1639_ = new_G1592_ & new_G1636_;
  assign new_G1648_ = new_G1596_ & new_G1645_;
  assign new_G1657_ = new_G1600_ & new_G1654_;
  assign new_G1666_ = new_G1604_ & new_G1663_;
  assign new_G1675_ = new_G1608_ & new_G1672_;
  assign new_G1895_ = new_G1893_ & new_G1894_;
  assign new_G1946_ = new_G1941_ | new_G1939_ | new_G1940_;
  assign new_G1998_ = new_G1996_ & new_G1997_;
  assign new_G2048_ = new_G2046_ & new_G2047_;
  assign new_G2103_ = new_G2101_ & new_G2102_;
  assign new_G2156_ = new_G2151_ | new_G2149_ | new_G2150_;
  assign new_G2210_ = new_G2208_ & new_G2209_;
  assign new_G2262_ = new_G2260_ & new_G2261_;
  assign new_G2271_ = ~new_G1892_;
  assign new_G2311_ = ~new_G2100_;
  assign new_G356_ = ~new_G619_ | ~new_G620_;
  assign new_G357_ = ~new_G582_ | ~new_G583_;
  assign new_G603_ = ~new_G3074_ | ~new_G3077_;
  assign new_G3078_ = ~new_G3074_;
  assign new_G606_ = ~new_G3066_ | ~new_G3069_;
  assign new_G3070_ = ~new_G3066_;
  assign new_G1670_ = new_G703_ & new_G1665_;
  assign new_G1679_ = new_G692_ & new_G1674_;
  assign new_G1942_ = new_G1933_ | new_G1936_;
  assign new_G1945_ = ~new_G1933_ & ~new_G1936_;
  assign new_G2152_ = new_G2143_ | new_G2146_;
  assign new_G2155_ = ~new_G2143_ & ~new_G2146_;
  assign new_G2445_ = new_G1993_ & new_G2293_;
  assign new_G2448_ = new_G2043_ & new_G2293_;
  assign new_G2455_ = new_G2205_ & new_G2302_;
  assign new_G2458_ = new_G2257_ & new_G2302_;
  assign new_G3142_ = new_G2328_;
  assign new_G3150_ = new_G2328_;
  assign new_G3208_ = new_G2375_;
  assign new_G3216_ = new_G2375_;
  assign G358 = ~new_G356_ | ~new_G357_;
  assign new_G604_ = ~new_G3071_ | ~new_G3078_;
  assign new_G607_ = ~new_G3063_ | ~new_G3070_;
  assign new_G1947_ = new_G1945_ & new_G1946_;
  assign new_G2157_ = new_G2155_ & new_G2156_;
  assign new_G2317_ = new_G1895_;
  assign new_G2338_ = new_G1998_;
  assign new_G2351_ = new_G2048_;
  assign new_G2364_ = new_G2103_;
  assign new_G2380_ = new_G2210_;
  assign new_G2388_ = new_G2262_;
  assign new_G605_ = ~new_G603_ | ~new_G604_;
  assign new_G608_ = ~new_G606_ | ~new_G607_;
  assign new_G2272_ = ~new_G1895_ | ~new_G1942_;
  assign new_G2312_ = ~new_G2103_ | ~new_G2152_;
  assign new_G3146_ = ~new_G3142_;
  assign new_G3154_ = ~new_G3150_;
  assign new_G3220_ = ~new_G3216_;
  assign new_G3212_ = ~new_G3208_;
  assign new_G2444_ = new_G1942_ & new_G2288_;
  assign new_G2451_ = new_G2448_;
  assign new_G2454_ = new_G2152_ & new_G2293_;
  assign new_G2461_ = new_G2458_;
  assign new_G2530_ = ~new_G2445_;
  assign new_G3323_ = new_G2458_;
  assign new_G349_ = ~new_G605_;
  assign new_G350_ = ~new_G608_;
  assign new_G2265_ = new_G2048_ & new_G1998_ & new_G1895_ & new_G1947_;
  assign new_G2273_ = ~new_G1993_ | ~new_G1895_ | ~new_G1947_;
  assign new_G2274_ = ~new_G1895_ | ~new_G1998_ | ~new_G2043_ | ~new_G1947_;
  assign new_G2309_ = new_G2262_ & new_G2210_ & new_G2103_ & new_G2157_;
  assign new_G2313_ = ~new_G2205_ | ~new_G2103_ | ~new_G2157_;
  assign new_G2314_ = ~new_G2103_ | ~new_G2210_ | ~new_G2257_ | ~new_G2157_;
  assign new_G2325_ = new_G1947_;
  assign new_G2372_ = new_G2157_;
  assign new_G2523_ = ~new_G2444_;
  assign new_G2533_ = ~new_G2454_;
  assign new_G3121_ = new_G2317_;
  assign new_G3131_ = new_G2317_;
  assign new_G3155_ = new_G2338_;
  assign new_G3163_ = new_G2338_;
  assign new_G3171_ = new_G2351_;
  assign new_G3179_ = new_G2351_;
  assign new_G3187_ = new_G2364_;
  assign new_G3197_ = new_G2364_;
  assign new_G3221_ = new_G2380_;
  assign new_G3229_ = new_G2380_;
  assign new_G3237_ = new_G2388_;
  assign new_G3245_ = new_G2388_;
  assign G351 = ~new_G349_ | ~new_G350_;
  assign new_G2275_ = ~new_G2274_ | ~new_G2273_ | ~new_G2271_ | ~new_G2272_;
  assign new_G2315_ = ~new_G2314_ | ~new_G2313_ | ~new_G2311_ | ~new_G2312_;
  assign new_G3329_ = ~new_G3323_;
  assign G372 = new_G2309_ & new_G2265_;
  assign new_G2324_ = ~new_G3131_ | ~new_G3138_;
  assign new_G2350_ = ~new_G3163_ | ~new_G3170_;
  assign new_G2363_ = ~new_G3179_ | ~new_G3186_;
  assign new_G2371_ = ~new_G3197_ | ~new_G3204_;
  assign new_G2387_ = ~new_G3229_ | ~new_G3236_;
  assign new_G2400_ = ~new_G3245_ | ~new_G3252_;
  assign new_G2268_ = new_G2265_;
  assign new_G3137_ = ~new_G3131_;
  assign new_G3161_ = ~new_G3155_;
  assign new_G2345_ = ~new_G3155_ | ~new_G3162_;
  assign new_G3169_ = ~new_G3163_;
  assign new_G3177_ = ~new_G3171_;
  assign new_G2358_ = ~new_G3171_ | ~new_G3178_;
  assign new_G3185_ = ~new_G3179_;
  assign new_G3203_ = ~new_G3197_;
  assign new_G3235_ = ~new_G3229_;
  assign new_G3243_ = ~new_G3237_;
  assign new_G2395_ = ~new_G3237_ | ~new_G3244_;
  assign new_G3251_ = ~new_G3245_;
  assign new_G3227_ = ~new_G3221_;
  assign new_G2432_ = ~new_G3221_ | ~new_G3228_;
  assign new_G2490_ = new_G2309_ & new_G2485_;
  assign new_G3127_ = ~new_G3121_;
  assign new_G3130_ = ~new_G3121_ | ~new_G3128_;
  assign new_G3139_ = new_G2325_;
  assign new_G3147_ = new_G2325_;
  assign new_G3193_ = ~new_G3187_;
  assign new_G3196_ = ~new_G3187_ | ~new_G3194_;
  assign new_G3205_ = new_G2372_;
  assign new_G3213_ = new_G2372_;
  assign new_G2307_ = ~new_G2265_ | ~new_G2315_;
  assign new_G2308_ = ~new_G2275_;
  assign new_G2323_ = ~new_G3134_ | ~new_G3137_;
  assign new_G2349_ = ~new_G3166_ | ~new_G3169_;
  assign new_G2362_ = ~new_G3182_ | ~new_G3185_;
  assign new_G2370_ = ~new_G3200_ | ~new_G3203_;
  assign new_G2386_ = ~new_G3232_ | ~new_G3235_;
  assign new_G2399_ = ~new_G3248_ | ~new_G3251_;
  assign new_G2344_ = ~new_G3158_ | ~new_G3161_;
  assign new_G2357_ = ~new_G3174_ | ~new_G3177_;
  assign new_G2394_ = ~new_G3240_ | ~new_G3243_;
  assign new_G2431_ = ~new_G3224_ | ~new_G3227_;
  assign new_G2464_ = new_G2315_ & new_G2302_;
  assign new_G2491_ = new_G2489_ | new_G2490_;
  assign new_G3129_ = ~new_G3124_ | ~new_G3127_;
  assign new_G3195_ = ~new_G3190_ | ~new_G3193_;
  assign new_G368_ = new_G2307_ & new_G2308_;
  assign new_G1615_ = ~new_G2323_ | ~new_G2324_;
  assign new_G2337_ = ~new_G3147_ | ~new_G3154_;
  assign new_G1633_ = ~new_G2349_ | ~new_G2350_;
  assign new_G1642_ = ~new_G2362_ | ~new_G2363_;
  assign new_G1651_ = ~new_G2370_ | ~new_G2371_;
  assign new_G2379_ = ~new_G3213_ | ~new_G3220_;
  assign new_G1669_ = ~new_G2386_ | ~new_G2387_;
  assign new_G1678_ = ~new_G2399_ | ~new_G2400_;
  assign new_G3145_ = ~new_G3139_;
  assign new_G2332_ = ~new_G3139_ | ~new_G3146_;
  assign new_G3153_ = ~new_G3147_;
  assign new_G2346_ = ~new_G2344_ | ~new_G2345_;
  assign new_G2359_ = ~new_G2357_ | ~new_G2358_;
  assign new_G3219_ = ~new_G3213_;
  assign new_G2396_ = ~new_G2394_ | ~new_G2395_;
  assign new_G3211_ = ~new_G3205_;
  assign new_G2425_ = ~new_G3205_ | ~new_G3212_;
  assign new_G2433_ = ~new_G2431_ | ~new_G2432_;
  assign new_G3272_ = ~new_G3129_ | ~new_G3130_;
  assign new_G3308_ = ~new_G3195_ | ~new_G3196_;
  assign G369 = ~new_G368_;
  assign new_G1613_ = ~new_G1615_;
  assign new_G2336_ = ~new_G3150_ | ~new_G3153_;
  assign new_G1631_ = ~new_G1633_;
  assign new_G1640_ = ~new_G1642_;
  assign new_G1649_ = ~new_G1651_;
  assign new_G2378_ = ~new_G3216_ | ~new_G3219_;
  assign new_G1667_ = ~new_G1669_;
  assign new_G1676_ = ~new_G1678_;
  assign new_G2331_ = ~new_G3142_ | ~new_G3145_;
  assign new_G2424_ = ~new_G3208_ | ~new_G3211_;
  assign new_G2467_ = new_G2464_;
  assign new_G2495_ = new_G2491_;
  assign new_G3295_ = new_G2464_;
  assign new_G3374_ = G330 & new_G2491_;
  assign new_G1614_ = new_G1613_ & new_G1610_;
  assign new_G1624_ = ~new_G2336_ | ~new_G2337_;
  assign new_G1632_ = new_G1631_ & new_G1628_;
  assign new_G1641_ = new_G1640_ & new_G1637_;
  assign new_G1650_ = new_G1649_ & new_G1646_;
  assign new_G1660_ = ~new_G2378_ | ~new_G2379_;
  assign new_G1668_ = new_G1667_ & new_G1664_;
  assign new_G1677_ = new_G1676_ & new_G1673_;
  assign new_G2333_ = ~new_G2331_ | ~new_G2332_;
  assign new_G2406_ = new_G2346_;
  assign new_G2409_ = new_G2346_;
  assign new_G2415_ = new_G2359_;
  assign new_G2419_ = new_G2359_;
  assign new_G2426_ = ~new_G2424_ | ~new_G2425_;
  assign new_G2439_ = new_G2396_;
  assign new_G2518_ = new_G2433_ & new_G2461_;
  assign new_G3276_ = ~new_G3272_;
  assign new_G3312_ = ~new_G3308_;
  assign new_G2612_ = G330 & new_G2396_;
  assign new_G3326_ = new_G2433_;
  assign new_G1617_ = ~new_G1616_ & ~new_G1612_ & ~new_G1614_;
  assign new_G1622_ = ~new_G1624_;
  assign new_G1635_ = ~new_G1634_ & ~new_G1630_ & ~new_G1632_;
  assign new_G1644_ = ~new_G1643_ & ~new_G1639_ & ~new_G1641_;
  assign new_G1653_ = ~new_G1652_ & ~new_G1648_ & ~new_G1650_;
  assign new_G1658_ = ~new_G1660_;
  assign new_G1671_ = ~new_G1670_ & ~new_G1666_ & ~new_G1668_;
  assign new_G1680_ = ~new_G1679_ & ~new_G1675_ & ~new_G1677_;
  assign new_G2500_ = new_G2467_ & new_G2268_;
  assign new_G2505_ = new_G2495_ & new_G2268_;
  assign new_G2519_ = new_G2455_ | new_G2518_;
  assign new_G3378_ = ~new_G3374_;
  assign new_G2642_ = ~new_G2467_;
  assign new_G2645_ = new_G2467_;
  assign new_G3301_ = ~new_G3295_;
  assign new_G1623_ = new_G1622_ & new_G1619_;
  assign new_G1659_ = new_G1658_ & new_G1655_;
  assign new_G2401_ = new_G2333_;
  assign new_G2501_ = new_G2275_ | new_G2500_;
  assign new_G2511_ = new_G2409_ & new_G2495_ & new_G2419_;
  assign new_G2512_ = new_G2495_ & new_G2415_;
  assign new_G2513_ = new_G2426_ & new_G2439_ & new_G2433_;
  assign new_G2514_ = new_G2439_ & new_G2433_;
  assign new_G2517_ = new_G2467_ & new_G2415_;
  assign new_G2531_ = ~new_G2409_ | ~new_G2451_;
  assign new_G2532_ = ~new_G2467_ | ~new_G2409_ | ~new_G2419_;
  assign new_G2534_ = ~new_G2426_ | ~new_G2455_;
  assign new_G2535_ = ~new_G2461_ | ~new_G2426_ | ~new_G2433_;
  assign new_G2607_ = ~new_G3326_ | ~new_G3329_;
  assign new_G3330_ = ~new_G3326_;
  assign new_G2643_ = new_G2642_ & G330 & new_G2491_;
  assign new_G2687_ = new_G1617_ & new_G2680_;
  assign new_G2725_ = new_G1635_ & new_G2718_;
  assign new_G2742_ = new_G1644_ & new_G2735_;
  assign new_G2760_ = new_G1653_ & new_G2753_;
  assign new_G2794_ = new_G1671_ & new_G2787_;
  assign new_G2811_ = new_G1680_ & new_G2804_;
  assign new_G3280_ = new_G2333_;
  assign new_G3290_ = new_G2409_;
  assign new_G3298_ = new_G2415_;
  assign new_G3316_ = new_G2426_;
  assign new_G3406_ = new_G2612_;
  assign new_G3414_ = new_G2612_;
  assign new_G3422_ = new_G2439_ & new_G2439_;
  assign new_G1626_ = ~new_G1625_ & ~new_G1621_ & ~new_G1623_;
  assign new_G1662_ = ~new_G1661_ & ~new_G1657_ & ~new_G1659_;
  assign new_G2567_ = G330 & new_G2512_;
  assign new_G2589_ = G330 & new_G2513_;
  assign new_G2608_ = ~new_G3323_ | ~new_G3330_;
  assign new_G2654_ = new_G2519_;
  assign new_G3253_ = new_G2505_;
  assign new_G3277_ = ~new_G2532_ | ~new_G2530_ | ~new_G2531_;
  assign new_G3287_ = new_G2448_ | new_G2517_;
  assign new_G3305_ = ~new_G2535_ | ~new_G2533_ | ~new_G2534_;
  assign new_G3313_ = new_G2519_;
  assign new_G3350_ = G330 & new_G2511_;
  assign new_G932_ = new_G2643_ | new_G2645_;
  assign new_G2508_ = new_G2419_ & new_G2409_ & new_G2495_ & new_G2401_;
  assign new_G2524_ = ~new_G2401_ | ~new_G2445_;
  assign new_G2525_ = ~new_G2451_ | ~new_G2401_ | ~new_G2406_;
  assign new_G2526_ = ~new_G2467_ | ~new_G2419_ | ~new_G2401_ | ~new_G2406_;
  assign new_G3294_ = ~new_G3290_;
  assign new_G2609_ = ~new_G2607_ | ~new_G2608_;
  assign new_G3410_ = ~new_G3406_;
  assign new_G3418_ = ~new_G3414_;
  assign new_G2624_ = ~new_G3422_ | ~new_G3425_;
  assign new_G3426_ = ~new_G3422_;
  assign new_G2629_ = new_G2501_;
  assign new_G2647_ = ~new_G2643_ & ~new_G2645_;
  assign new_G2706_ = new_G1626_ & new_G2699_;
  assign new_G2777_ = new_G1662_ & new_G2770_;
  assign new_G3264_ = new_G2501_;
  assign new_G3284_ = ~new_G3280_;
  assign new_G3302_ = ~new_G3298_;
  assign new_G3303_ = ~new_G3298_ | ~new_G3301_;
  assign new_G3320_ = ~new_G3316_;
  assign new_G3398_ = G330 & new_G2514_;
  assign new_G2657_ = ~new_G2654_;
  assign new_G398_ = new_G2519_ & new_G2654_;
  assign new_G933_ = new_G932_ & new_G927_;
  assign new_G2527_ = ~new_G2526_ | ~new_G2525_ | ~new_G2523_ | ~new_G2524_;
  assign new_G3259_ = ~new_G3253_;
  assign new_G3354_ = ~new_G3350_;
  assign new_G3293_ = ~new_G3287_;
  assign new_G2563_ = ~new_G3287_ | ~new_G3294_;
  assign new_G3311_ = ~new_G3305_;
  assign new_G2585_ = ~new_G3305_ | ~new_G3312_;
  assign new_G2625_ = ~new_G3419_ | ~new_G3426_;
  assign new_G3283_ = ~new_G3277_;
  assign new_G3286_ = ~new_G3277_ | ~new_G3284_;
  assign new_G3304_ = ~new_G3295_ | ~new_G3302_;
  assign new_G3319_ = ~new_G3313_;
  assign new_G3322_ = ~new_G3313_ | ~new_G3320_;
  assign new_G3358_ = new_G2567_;
  assign new_G3366_ = new_G2567_;
  assign new_G3382_ = new_G2589_;
  assign new_G3390_ = new_G2589_;
  assign new_G397_ = new_G2657_ & G330 & new_G2514_;
  assign new_G2544_ = G330 & new_G2508_;
  assign new_G2562_ = ~new_G3290_ | ~new_G3293_;
  assign new_G2584_ = ~new_G3308_ | ~new_G3311_;
  assign new_G3402_ = ~new_G3398_;
  assign new_G2626_ = ~new_G2624_ | ~new_G2625_;
  assign new_G2632_ = ~new_G2629_;
  assign new_G2634_ = new_G2501_ & new_G2629_;
  assign new_G2650_ = new_G2647_;
  assign new_G3268_ = ~new_G3264_;
  assign new_G3256_ = new_G2508_;
  assign new_G3285_ = ~new_G3280_ | ~new_G3283_;
  assign new_G3321_ = ~new_G3316_ | ~new_G3319_;
  assign new_G3371_ = ~new_G3303_ | ~new_G3304_;
  assign new_G3403_ = new_G2609_;
  assign new_G3411_ = new_G2609_;
  assign new_G362_ = new_G938_ | new_G929_ | new_G933_;
  assign new_G1030_ = ~new_G938_ & ~new_G929_ & ~new_G933_;
  assign G399 = new_G397_ | new_G398_;
  assign new_G2564_ = ~new_G2562_ | ~new_G2563_;
  assign new_G3362_ = ~new_G3358_;
  assign new_G3370_ = ~new_G3366_;
  assign new_G2586_ = ~new_G2584_ | ~new_G2585_;
  assign new_G3386_ = ~new_G3382_;
  assign new_G3394_ = ~new_G3390_;
  assign new_G2633_ = new_G2632_ & G330 & new_G2505_;
  assign new_G3261_ = new_G2527_;
  assign new_G3269_ = new_G2527_;
  assign new_G3347_ = ~new_G3285_ | ~new_G3286_;
  assign new_G3395_ = ~new_G3321_ | ~new_G3322_;
  assign new_G363_ = ~new_G1030_;
  assign new_G2536_ = ~new_G3256_ | ~new_G3259_;
  assign new_G3260_ = ~new_G3256_;
  assign new_G3377_ = ~new_G3371_;
  assign new_G2580_ = ~new_G3371_ | ~new_G3378_;
  assign new_G3409_ = ~new_G3403_;
  assign new_G2616_ = ~new_G3403_ | ~new_G3410_;
  assign new_G3417_ = ~new_G3411_;
  assign new_G2622_ = ~new_G3411_ | ~new_G3418_;
  assign new_G2635_ = ~new_G2633_ & ~new_G2634_;
  assign new_G2805_ = new_G2626_ & new_G2802_;
  assign new_G2808_ = new_G2626_ & new_G2803_;
  assign new_G3334_ = new_G2544_;
  assign new_G3342_ = new_G2544_;
  assign new_G3454_ = new_G2650_;
  assign G364 = new_G362_ & new_G363_;
  assign new_G2537_ = ~new_G3253_ | ~new_G3260_;
  assign new_G3275_ = ~new_G3269_;
  assign new_G2540_ = ~new_G3269_ | ~new_G3276_;
  assign new_G3353_ = ~new_G3347_;
  assign new_G2557_ = ~new_G3347_ | ~new_G3354_;
  assign new_G2579_ = ~new_G3374_ | ~new_G3377_;
  assign new_G3401_ = ~new_G3395_;
  assign new_G2602_ = ~new_G3395_ | ~new_G3402_;
  assign new_G2615_ = ~new_G3406_ | ~new_G3409_;
  assign new_G2621_ = ~new_G3414_ | ~new_G3417_;
  assign new_G3267_ = ~new_G3261_;
  assign new_G3112_ = ~new_G3261_ | ~new_G3268_;
  assign new_G3355_ = new_G2564_;
  assign new_G3363_ = new_G2564_;
  assign new_G3379_ = new_G2586_;
  assign new_G3387_ = new_G2586_;
  assign new_G2538_ = ~new_G2536_ | ~new_G2537_;
  assign new_G2539_ = ~new_G3272_ | ~new_G3275_;
  assign new_G3338_ = ~new_G3334_;
  assign new_G3346_ = ~new_G3342_;
  assign new_G2556_ = ~new_G3350_ | ~new_G3353_;
  assign new_G2581_ = ~new_G2579_ | ~new_G2580_;
  assign new_G2601_ = ~new_G3398_ | ~new_G3401_;
  assign new_G2617_ = ~new_G2615_ | ~new_G2616_;
  assign new_G2623_ = ~new_G2621_ | ~new_G2622_;
  assign new_G2638_ = new_G2635_;
  assign new_G3458_ = ~new_G3454_;
  assign new_G2814_ = new_G2811_ | new_G2805_ | new_G2808_;
  assign new_G2816_ = ~new_G2811_ & ~new_G2805_ & ~new_G2808_;
  assign new_G3111_ = ~new_G3264_ | ~new_G3267_;
  assign new_G2541_ = ~new_G2539_ | ~new_G2540_;
  assign new_G2558_ = ~new_G2556_ | ~new_G2557_;
  assign new_G3361_ = ~new_G3355_;
  assign new_G2571_ = ~new_G3355_ | ~new_G3362_;
  assign new_G3369_ = ~new_G3363_;
  assign new_G2577_ = ~new_G3363_ | ~new_G3370_;
  assign new_G3385_ = ~new_G3379_;
  assign new_G2593_ = ~new_G3379_ | ~new_G3386_;
  assign new_G3393_ = ~new_G3387_;
  assign new_G2598_ = ~new_G3387_ | ~new_G3394_;
  assign new_G2603_ = ~new_G2601_ | ~new_G2602_;
  assign new_G3113_ = ~new_G3111_ | ~new_G3112_;
  assign new_G3116_ = G330 & new_G2538_;
  assign new_G3451_ = ~new_G2623_;
  assign new_G395_ = ~new_G2816_;
  assign new_G2570_ = ~new_G3358_ | ~new_G3361_;
  assign new_G2576_ = ~new_G3366_ | ~new_G3369_;
  assign new_G2592_ = ~new_G3382_ | ~new_G3385_;
  assign new_G2597_ = ~new_G3390_ | ~new_G3393_;
  assign new_G2736_ = new_G2581_ & new_G2733_;
  assign new_G2739_ = new_G2581_ & new_G2734_;
  assign new_G2788_ = new_G2617_ & new_G2785_;
  assign new_G3438_ = new_G2638_;
  assign new_G3446_ = new_G2617_ & new_G2647_;
  assign new_G3459_ = new_G2814_;
  assign G396 = new_G2814_ & new_G395_;
  assign new_G3119_ = ~new_G3113_;
  assign new_G3120_ = ~new_G3116_;
  assign new_G2572_ = ~new_G2570_ | ~new_G2571_;
  assign new_G2578_ = ~new_G2576_ | ~new_G2577_;
  assign new_G2594_ = ~new_G2592_ | ~new_G2593_;
  assign new_G2599_ = ~new_G2597_ | ~new_G2598_;
  assign new_G2677_ = ~new_G3451_ | ~new_G3458_;
  assign new_G3457_ = ~new_G3451_;
  assign new_G2700_ = new_G2558_ & new_G2697_;
  assign new_G2771_ = new_G2603_ & new_G2768_;
  assign new_G3331_ = new_G2541_;
  assign new_G3339_ = new_G2541_;
  assign new_G3427_ = new_G2558_;
  assign new_G3443_ = new_G2603_;
  assign new_G954_ = ~new_G3116_ | ~new_G3119_;
  assign new_G955_ = ~new_G3113_ | ~new_G3120_;
  assign new_G2600_ = ~new_G2599_;
  assign new_G3442_ = ~new_G3438_;
  assign new_G3450_ = ~new_G3446_;
  assign new_G2676_ = ~new_G3454_ | ~new_G3457_;
  assign new_G2745_ = new_G2742_ | new_G2736_ | new_G2739_;
  assign new_G2748_ = ~new_G2742_ & ~new_G2736_ & ~new_G2739_;
  assign new_G3465_ = ~new_G3459_;
  assign new_G3435_ = ~new_G2578_;
  assign new_G950_ = ~new_G954_ | ~new_G955_;
  assign new_G3337_ = ~new_G3331_;
  assign new_G2548_ = ~new_G3331_ | ~new_G3338_;
  assign new_G3345_ = ~new_G3339_;
  assign new_G2553_ = ~new_G3339_ | ~new_G3346_;
  assign new_G2661_ = ~new_G2600_ & ~new_G2650_;
  assign new_G2662_ = new_G2650_ & new_G2594_ & new_G2617_ & new_G2603_;
  assign new_G3433_ = ~new_G3427_;
  assign new_G3449_ = ~new_G3443_;
  assign new_G2672_ = ~new_G3443_ | ~new_G3450_;
  assign new_G2674_ = ~new_G2676_ | ~new_G2677_;
  assign new_G2719_ = new_G2572_ & new_G2716_;
  assign new_G2754_ = new_G2594_ & new_G2751_;
  assign new_G3430_ = new_G2572_ & new_G2635_;
  assign new_G383_ = ~new_G2748_;
  assign new_G951_ = new_G950_ & new_G943_;
  assign new_G2547_ = ~new_G3334_ | ~new_G3337_;
  assign new_G2552_ = ~new_G3342_ | ~new_G3345_;
  assign new_G2663_ = new_G2661_ | new_G2662_;
  assign new_G2670_ = ~new_G3435_ | ~new_G3442_;
  assign new_G3441_ = ~new_G3435_;
  assign new_G2671_ = ~new_G3446_ | ~new_G3449_;
  assign new_G2675_ = ~new_G2674_;
  assign new_G3491_ = new_G2745_;
  assign new_G3499_ = new_G2745_;
  assign G384 = new_G2745_ & new_G383_;
  assign new_G2549_ = ~new_G2547_ | ~new_G2548_;
  assign new_G2554_ = ~new_G2552_ | ~new_G2553_;
  assign new_G2664_ = ~new_G3430_ | ~new_G3433_;
  assign new_G3434_ = ~new_G3430_;
  assign new_G2669_ = ~new_G3438_ | ~new_G3441_;
  assign new_G2673_ = ~new_G2671_ | ~new_G2672_;
  assign new_G2757_ = new_G2663_ & new_G2752_;
  assign new_G2791_ = new_G2675_ & new_G2786_;
  assign new_G365_ = new_G951_ | new_G944_ | new_G947_;
  assign new_G1031_ = ~new_G951_ & ~new_G944_ & ~new_G947_;
  assign new_G2555_ = ~new_G2554_;
  assign new_G2665_ = ~new_G3427_ | ~new_G3434_;
  assign new_G2667_ = ~new_G2669_ | ~new_G2670_;
  assign new_G2774_ = new_G2673_ & new_G2769_;
  assign new_G3497_ = ~new_G3491_;
  assign new_G3505_ = ~new_G3499_;
  assign new_G366_ = ~new_G1031_;
  assign new_G2658_ = ~new_G2555_ & ~new_G2638_;
  assign new_G2659_ = new_G2638_ & new_G2549_ & new_G2572_ & new_G2558_;
  assign new_G2666_ = ~new_G2664_ | ~new_G2665_;
  assign new_G2668_ = ~new_G2667_;
  assign new_G2681_ = new_G2549_ & new_G2678_;
  assign new_G2763_ = new_G2760_ | new_G2754_ | new_G2757_;
  assign new_G2765_ = ~new_G2760_ & ~new_G2754_ & ~new_G2757_;
  assign new_G2797_ = new_G2794_ | new_G2788_ | new_G2791_;
  assign new_G2799_ = ~new_G2794_ & ~new_G2788_ & ~new_G2791_;
  assign G367 = new_G365_ & new_G366_;
  assign new_G2660_ = new_G2658_ | new_G2659_;
  assign new_G2703_ = new_G2666_ & new_G2698_;
  assign new_G2722_ = new_G2668_ & new_G2717_;
  assign new_G2780_ = new_G2777_ | new_G2771_ | new_G2774_;
  assign new_G2782_ = ~new_G2777_ & ~new_G2771_ & ~new_G2774_;
  assign new_G386_ = ~new_G2765_;
  assign new_G392_ = ~new_G2799_;
  assign new_G2684_ = new_G2660_ & new_G2679_;
  assign new_G3462_ = new_G2797_;
  assign new_G3470_ = new_G2763_;
  assign G387 = new_G2763_ & new_G386_;
  assign new_G389_ = ~new_G2782_;
  assign G393 = new_G2797_ & new_G392_;
  assign new_G2709_ = new_G2706_ | new_G2700_ | new_G2703_;
  assign new_G2713_ = ~new_G2706_ & ~new_G2700_ & ~new_G2703_;
  assign new_G2728_ = new_G2725_ | new_G2719_ | new_G2722_;
  assign new_G2730_ = ~new_G2725_ & ~new_G2719_ & ~new_G2722_;
  assign new_G2922_ = new_G2765_ & new_G2782_ & new_G2816_ & new_G2799_;
  assign new_G3467_ = new_G2780_;
  assign G390 = new_G2780_ & new_G389_;
  assign new_G2690_ = new_G2687_ | new_G2681_ | new_G2684_;
  assign new_G2694_ = ~new_G2687_ & ~new_G2681_ & ~new_G2684_;
  assign new_G2821_ = ~new_G3462_ | ~new_G3465_;
  assign new_G3466_ = ~new_G3462_;
  assign new_G3474_ = ~new_G3470_;
  assign G378 = new_G2709_ & new_G2709_;
  assign new_G380_ = ~new_G2730_;
  assign new_G2822_ = ~new_G3459_ | ~new_G3466_;
  assign new_G3473_ = ~new_G3467_;
  assign new_G2827_ = ~new_G3467_ | ~new_G3474_;
  assign new_G2839_ = new_G2728_;
  assign new_G2883_ = new_G2709_ & new_G2871_;
  assign new_G3507_ = new_G2709_;
  assign G375 = new_G2690_ & new_G2690_;
  assign G381 = new_G2728_ & new_G380_;
  assign new_G2823_ = ~new_G2821_ | ~new_G2822_;
  assign new_G2826_ = ~new_G3470_ | ~new_G3473_;
  assign new_G2880_ = new_G2871_ & new_G2690_;
  assign new_G2925_ = new_G2694_ & new_G2713_ & new_G2748_ & new_G2730_;
  assign new_G2928_ = new_G2874_ & new_G2713_ & new_G2694_;
  assign new_G3510_ = new_G2690_;
  assign new_G2828_ = ~new_G2826_ | ~new_G2827_;
  assign new_G3494_ = new_G2839_;
  assign new_G3502_ = new_G2839_;
  assign new_G3513_ = ~new_G3507_;
  assign new_G3544_ = new_G2883_;
  assign new_G3552_ = new_G2883_;
  assign new_G406_ = new_G2922_ & new_G2925_;
  assign new_G2929_ = new_G2922_ & new_G2925_;
  assign new_G3475_ = new_G2823_;
  assign new_G3483_ = new_G2823_;
  assign new_G3514_ = ~new_G3510_;
  assign new_G3515_ = ~new_G3510_ | ~new_G3513_;
  assign new_G3541_ = new_G2880_;
  assign new_G3549_ = new_G2880_;
  assign G407 = ~new_G406_;
  assign new_G2930_ = ~new_G2928_ & ~new_G2929_;
  assign new_G2842_ = ~new_G3494_ | ~new_G3497_;
  assign new_G3498_ = ~new_G3494_;
  assign new_G2852_ = ~new_G3502_ | ~new_G3505_;
  assign new_G3506_ = ~new_G3502_;
  assign new_G3548_ = ~new_G3544_;
  assign new_G3556_ = ~new_G3552_;
  assign new_G3478_ = new_G2828_;
  assign new_G3486_ = new_G2828_;
  assign new_G3516_ = ~new_G3507_ | ~new_G3514_;
  assign new_G408_ = G213 & new_G2930_;
  assign new_G3481_ = ~new_G3475_;
  assign new_G3489_ = ~new_G3483_;
  assign new_G2843_ = ~new_G3491_ | ~new_G3498_;
  assign new_G2853_ = ~new_G3499_ | ~new_G3506_;
  assign new_G3547_ = ~new_G3541_;
  assign new_G2887_ = ~new_G3541_ | ~new_G3548_;
  assign new_G2896_ = ~new_G3549_ | ~new_G3556_;
  assign new_G3555_ = ~new_G3549_;
  assign new_G3520_ = ~new_G3515_ | ~new_G3516_;
  assign G409 = ~new_G408_;
  assign new_G2831_ = ~new_G3478_ | ~new_G3481_;
  assign new_G3482_ = ~new_G3478_;
  assign new_G2836_ = ~new_G3486_ | ~new_G3489_;
  assign new_G3490_ = ~new_G3486_;
  assign new_G2844_ = ~new_G2842_ | ~new_G2843_;
  assign new_G2848_ = ~new_G2852_ | ~new_G2853_;
  assign new_G2886_ = ~new_G3544_ | ~new_G3547_;
  assign new_G2895_ = ~new_G3552_ | ~new_G3555_;
  assign new_G2832_ = ~new_G3475_ | ~new_G3482_;
  assign new_G2837_ = ~new_G3483_ | ~new_G3490_;
  assign new_G2849_ = ~new_G2848_;
  assign new_G3524_ = ~new_G3520_;
  assign new_G2888_ = ~new_G2886_ | ~new_G2887_;
  assign new_G2891_ = ~new_G2895_ | ~new_G2896_;
  assign new_G2833_ = ~new_G2831_ | ~new_G2832_;
  assign new_G2838_ = ~new_G2836_ | ~new_G2837_;
  assign new_G2892_ = ~new_G2891_;
  assign new_G3517_ = new_G2844_;
  assign new_G2906_ = new_G2900_ & new_G2844_ & new_G2888_;
  assign new_G2908_ = new_G2903_ & new_G2849_ & new_G2888_;
  assign new_G2913_ = ~new_G2838_;
  assign new_G3523_ = ~new_G3517_;
  assign new_G2855_ = ~new_G3517_ | ~new_G3524_;
  assign new_G2907_ = new_G2903_ & new_G2844_ & new_G2892_;
  assign new_G2909_ = new_G2900_ & new_G2849_ & new_G2892_;
  assign new_G3525_ = new_G2833_;
  assign new_G3533_ = new_G2833_;
  assign new_G2854_ = ~new_G3520_ | ~new_G3523_;
  assign new_G2910_ = new_G2909_ | new_G2908_ | new_G2906_ | new_G2907_;
  assign new_G3560_ = new_G2913_;
  assign new_G3568_ = new_G2913_;
  assign new_G2856_ = ~new_G2854_ | ~new_G2855_;
  assign new_G3539_ = ~new_G3533_;
  assign new_G3531_ = ~new_G3525_;
  assign new_G3572_ = ~new_G3568_;
  assign new_G3564_ = ~new_G3560_;
  assign new_G3557_ = new_G2910_;
  assign new_G3565_ = new_G2910_;
  assign new_G3528_ = new_G2856_;
  assign new_G3536_ = new_G2856_;
  assign new_G2921_ = ~new_G3557_ | ~new_G3564_;
  assign new_G2917_ = ~new_G3565_ | ~new_G3572_;
  assign new_G3571_ = ~new_G3565_;
  assign new_G3563_ = ~new_G3557_;
  assign new_G2863_ = ~new_G3528_ | ~new_G3531_;
  assign new_G2859_ = ~new_G3536_ | ~new_G3539_;
  assign new_G2920_ = ~new_G3560_ | ~new_G3563_;
  assign new_G2916_ = ~new_G3568_ | ~new_G3571_;
  assign new_G3540_ = ~new_G3536_;
  assign new_G3532_ = ~new_G3528_;
  assign new_G2864_ = ~new_G3525_ | ~new_G3532_;
  assign new_G2860_ = ~new_G3533_ | ~new_G3540_;
  assign new_G403_ = ~new_G2920_ | ~new_G2921_;
  assign new_G404_ = ~new_G2916_ | ~new_G2917_;
  assign new_G400_ = ~new_G2863_ | ~new_G2864_;
  assign new_G401_ = ~new_G2859_ | ~new_G2860_;
  assign G405 = new_G403_ & new_G404_;
  assign G402 = ~new_G400_ | ~new_G401_;
endmodule


