// NOR_NOT mapped module c432

module c432 (
  input  G1gat   ,
  input  G4gat   ,
  input  G8gat   ,
  input  G11gat  ,
  input  G14gat  ,
  input  G17gat  ,
  input  G21gat  ,
  input  G24gat  ,
  input  G27gat  ,
  input  G30gat  ,
  input  G34gat  ,
  input  G37gat  ,
  input  G40gat  ,
  input  G43gat  ,
  input  G47gat  ,
  input  G50gat  ,
  input  G53gat  ,
  input  G56gat  ,
  input  G60gat  ,
  input  G63gat  ,
  input  G66gat  ,
  input  G69gat  ,
  input  G73gat  ,
  input  G76gat  ,
  input  G79gat  ,
  input  G82gat  ,
  input  G86gat  ,
  input  G89gat  ,
  input  G92gat  ,
  input  G95gat  ,
  input  G99gat  ,
  input  G102gat ,
  input  G105gat ,
  input  G108gat ,
  input  G112gat ,
  input  G115gat ,
  output G223gat ,
  output G329gat ,
  output G370gat ,
  output G421gat ,
  output G430gat ,
  output G431gat ,
  output G432gat );

  wire wr_8;
  wire wr_9;
  wire wr_10;
  wire wr_11;
  wire wr_12;
  wire wr_13;
  wire wr_14;
  wire wr_15;
  wire wr_16;
  wire wr_17;
  wire wr_18;
  wire wr_19;
  wire wr_20;
  wire wr_21;
  wire wr_22;
  wire wr_23;
  wire wr_24;
  wire wr_25;
  wire wr_26;
  wire wr_27;
  wire wr_28;
  wire wr_29;
  wire wr_30;
  wire wr_31;
  wire wr_32;
  wire wr_33;
  wire wr_34;
  wire wr_35;
  wire wr_36;
  wire wr_37;
  wire wr_38;
  wire wr_39;
  wire wr_40;
  wire wr_41;
  wire wr_42;
  wire wr_43;
  wire wr_44;
  wire wr_45;
  wire wr_46;
  wire wr_47;
  wire wr_48;
  wire wr_49;
  wire wr_50;
  wire wr_51;
  wire wr_52;
  wire wr_53;
  wire wr_54;
  wire wr_55;
  wire wr_56;
  wire wr_57;
  wire wr_58;
  wire wr_59;
  wire wr_60;
  wire wr_61;
  wire wr_62;
  wire wr_63;
  wire wr_64;
  wire wr_65;
  wire wr_66;
  wire wr_67;
  wire wr_68;
  wire wr_69;
  wire wr_70;
  wire wr_71;
  wire wr_72;
  wire wr_73;
  wire wr_74;
  wire wr_75;
  wire wr_76;
  wire wr_77;
  wire wr_78;
  wire wr_79;
  wire wr_80;
  wire wr_81;
  wire wr_82;
  wire wr_83;
  wire wr_84;
  wire wr_85;
  wire wr_86;
  wire wr_87;
  wire wr_88;
  wire wr_89;
  wire wr_90;
  wire wr_91;
  wire wr_92;
  wire wr_93;
  wire wr_94;
  wire wr_95;
  wire wr_96;
  wire wr_97;
  wire wr_98;
  wire wr_99;
  wire wr_100;
  wire wr_101;
  wire wr_102;
  wire wr_103;
  wire wr_104;
  wire wr_105;
  wire wr_106;
  wire wr_107;
  wire wr_108;
  wire wr_109;
  wire wr_110;
  wire wr_111;
  wire wr_112;
  wire wr_113;
  wire wr_114;
  wire wr_115;
  wire wr_116;
  wire wr_117;
  wire wr_118;
  wire wr_119;
  wire wr_120;
  wire wr_121;
  wire wr_122;
  wire wr_123;
  wire wr_124;
  wire wr_125;
  wire wr_126;
  wire wr_127;
  wire wr_128;
  wire wr_129;
  wire wr_130;
  wire wr_131;
  wire wr_132;
  wire wr_133;
  wire wr_134;
  wire wr_135;
  wire wr_136;
  wire wr_137;
  wire wr_138;
  wire wr_139;
  wire wr_140;
  wire wr_141;
  wire wr_142;
  wire wr_143;
  wire wr_144;
  wire wr_145;
  wire wr_146;
  wire wr_147;
  wire wr_148;
  wire wr_149;
  wire wr_150;
  wire wr_151;
  wire wr_152;
  wire wr_153;
  wire wr_154;
  wire wr_155;
  wire wr_156;
  wire wr_157;
  wire wr_158;
  wire wr_159;
  wire wr_160;
  wire wr_161;
  wire wr_162;
  wire wr_163;
  wire wr_164;
  wire wr_165;
  wire wr_166;
  wire wr_167;
  wire wr_168;
  wire wr_169;
  wire wr_170;
  wire wr_171;
  wire wr_172;
  wire wr_173;
  wire wr_174;
  wire wr_175;
  wire wr_176;
  wire wr_177;
  wire wr_178;
  wire wr_179;
  wire wr_180;
  wire wr_181;
  wire wr_182;
  wire wr_183;
  wire wr_184;
  wire wr_185;
  wire wr_186;
  wire wr_187;
  wire wr_188;
  wire wr_189;
  wire wr_190;
  wire wr_191;
  wire wr_192;
  wire wr_193;
  wire wr_194;
  wire wr_195;
  wire wr_196;
  wire wr_197;
  wire wr_198;
  wire wr_199;
  wire wr_200;
  wire wr_201;
  wire wr_202;
  wire wr_203;
  wire wr_204;
  wire wr_205;
  wire wr_206;
  wire wr_207;
  wire wr_208;
  wire wr_209;
  wire wr_210;
  wire wr_211;
  wire wr_212;
  wire wr_213;
  wire wr_214;
  wire wr_215;
  wire wr_216;
  wire wr_217;
  wire wr_218;
  wire wr_219;
  wire wr_220;
  wire wr_221;
  wire wr_222;
  wire wr_223;
  wire wr_224;
  wire wr_225;
  wire wr_226;
  wire wr_227;
  wire wr_228;
  wire wr_229;
  wire wr_230;
  wire wr_231;
  wire wr_232;
  wire wr_233;
  wire wr_234;
  wire wr_235;
  wire wr_236;
  wire wr_237;
  wire wr_238;
  wire wr_239;
  wire wr_240;
  wire wr_241;
  wire wr_242;
  wire wr_243;
  wire wr_244;
  wire wr_245;
  wire wr_246;
  wire wr_247;
  wire wr_248;
  wire wr_249;
  wire wr_250;
  wire wr_251;
  wire wr_252;
  wire wr_253;
  wire wr_254;
  wire wr_255;
  wire wr_256;
  wire wr_257;
  wire wr_258;
  wire wr_259;
  wire wr_260;
  wire wr_261;
  wire wr_262;
  wire wr_263;
  wire wr_264;
  wire wr_265;
  wire wr_266;
  wire wr_267;
  wire wr_268;
  wire wr_269;
  wire wr_270;
  wire wr_271;
  wire wr_272;
  wire wr_273;
  wire wr_274;
  wire wr_275;
  wire wr_276;
  wire wr_277;
  wire wr_278;
  wire wr_279;
  wire wr_280;
  wire wr_281;
  wire wr_282;
  wire wr_283;
  wire wr_284;
  wire wr_285;
  wire wr_286;
  wire wr_287;
  wire wr_288;
  wire wr_289;
  wire wr_290;
  wire wr_291;
  wire wr_292;
  wire wr_293;
  wire wr_294;
  wire wr_295;
  wire wr_296;
  wire wr_297;
  wire wr_298;
  wire wr_299;
  wire wr_300;
  wire wr_301;
  wire wr_302;
  wire wr_303;
  wire wr_304;
  wire wr_305;
  wire wr_306;
  wire wr_307;
  wire wr_308;
  wire wr_309;
  wire wr_310;
  wire wr_311;
  wire wr_312;
  wire wr_313;
  wire wr_314;
  wire wr_315;
  wire wr_316;
  wire wr_317;
  wire wr_318;
  wire wr_319;
  wire wr_320;
  wire wr_321;
  wire wr_322;
  wire wr_323;
  wire wr_324;
  wire wr_325;
  wire wr_326;
  wire wr_327;
  wire wr_328;
  wire wr_329;
  wire wr_330;
  wire wr_331;
  wire wr_332;
  wire wr_333;
  wire wr_334;
  wire wr_335;
  wire wr_336;
  wire wr_337;
  wire wr_338;
  wire wr_339;
  wire wr_340;
  wire wr_341;
  wire wr_342;
  wire wr_343;
  wire wr_344;
  wire wr_345;
  wire wr_346;
  wire wr_347;
  wire wr_348;
  wire wr_349;
  wire wr_350;
  wire wr_351;

  not    g1( wr_8    ,           G17gat  );
  not    g2( wr_10   ,           G4gat   );
  not    g3( wr_12   ,           G30gat  );
  not    g4( wr_14   ,           G43gat  );
  not    g5( wr_16   ,           G56gat  );
  not    g6( wr_18   ,           G69gat  );
  not    g7( wr_20   ,           G82gat  );
  not    g8( wr_22   ,           G108gat );
  not    g9( wr_24   ,           G95gat  );
  not   g10( wr_288  ,           G115gat );
  not   g11( wr_299  ,           G105gat );
  not   g12( wr_266  ,           G79gat  );
  not   g13( wr_277  ,           G92gat  );
  not   g14( wr_286  ,           G102gat );
  not   g15( wr_297  ,           G89gat  );
  not   g16( wr_255  ,           G66gat  );
  not   g17( wr_264  ,           G63gat  );
  not   g18( wr_275  ,           G76gat  );
  not   g19( wr_284  ,           G112gat );
  not   g20( wr_295  ,           G99gat  );
  not   g21( wr_222  ,           G40gat  );
  not   g22( wr_253  ,           G50gat  );
  not   g23( wr_244  ,           G53gat  );
  not   g24( wr_262  ,           G73gat  );
  not   g25( wr_273  ,           G86gat  );
  not   g26( wr_220  ,           G24gat  );
  not   g27( wr_251  ,           G60gat  );
  not   g28( wr_242  ,           G37gat  );
  not   g29( wr_218  ,           G34gat  );
  not   g30( wr_233  ,           G27gat  );
  not   g31( wr_240  ,           G47gat  );
  not   g32( wr_231  ,           G11gat  );
  not   g33( wr_209  ,           G14gat  );
  not   g34( wr_211  ,           G8gat   );
  not   g35( wr_229  ,           G21gat  );
  not   g36( wr_207  ,           G1gat   );
  nor   g37( wr_9    , wr_8    , G11gat  );
  nor   g38( wr_11   , wr_10   , G1gat   );
  nor   g39( wr_13   , wr_12   , G24gat  );
  nor   g40( wr_15   , wr_14   , G37gat  );
  nor   g41( wr_17   , wr_16   , G50gat  );
  nor   g42( wr_19   , wr_18   , G63gat  );
  nor   g43( wr_21   , wr_20   , G76gat  );
  nor   g44( wr_23   , wr_22   , G102gat );
  nor   g45( wr_25   , wr_24   , G89gat  );
  nor   g46( wr_42   , G21gat  , wr_8    );
  nor   g47( wr_46   , wr_10   , G1gat   );
  nor   g48( wr_48   , G8gat   , wr_10   );
  nor   g49( wr_52   , wr_12   , G24gat  );
  nor   g50( wr_54   , G34gat  , wr_12   );
  nor   g51( wr_61   , G47gat  , wr_14   );
  nor   g52( wr_68   , G60gat  , wr_16   );
  nor   g53( wr_75   , G73gat  , wr_18   );
  nor   g54( wr_82   , G86gat  , wr_20   );
  nor   g55( wr_89   , G112gat , wr_22   );
  nor   g56( wr_96   , G99gat  , wr_24   );
  nor   g57( wr_151  , G66gat  , wr_16   );
  nor   g58( wr_160  , G79gat  , wr_18   );
  nor   g59( wr_169  , G92gat  , wr_20   );
  nor   g60( wr_133  , G40gat  , wr_12   );
  nor   g61( wr_142  , G53gat  , wr_14   );
  nor   g62( wr_178  , G115gat , wr_22   );
  nor   g63( wr_187  , G105gat , wr_24   );
  nor   g64( wr_124  , G14gat  , wr_10   );
  nor   g65( wr_115  , G27gat  , wr_8    );
  nor   g66( wr_26   , wr_25   , wr_23   );
  not   g67( wr_43   ,           wr_42   );
  not   g68( wr_49   ,           wr_48   );
  not   g69( wr_55   ,           wr_54   );
  not   g70( wr_58   ,           wr_15   );
  not   g71( wr_62   ,           wr_61   );
  not   g72( wr_65   ,           wr_17   );
  not   g73( wr_69   ,           wr_68   );
  not   g74( wr_72   ,           wr_19   );
  not   g75( wr_76   ,           wr_75   );
  not   g76( wr_79   ,           wr_21   );
  not   g77( wr_83   ,           wr_82   );
  not   g78( wr_86   ,           wr_23   );
  not   g79( wr_90   ,           wr_89   );
  not   g80( wr_93   ,           wr_25   );
  not   g81( wr_97   ,           wr_96   );
  not   g82( wr_143  ,           wr_142  );
  not   g83( wr_152  ,           wr_151  );
  not   g84( wr_161  ,           wr_160  );
  not   g85( wr_170  ,           wr_169  );
  not   g86( wr_179  ,           wr_178  );
  not   g87( wr_188  ,           wr_187  );
  not   g88( wr_134  ,           wr_133  );
  not   g89( wr_125  ,           wr_124  );
  not   g90( wr_116  ,           wr_115  );
  not   g91( wr_27   ,           wr_26   );
  nor   g92( wr_28   , wr_27   , wr_21   );
  not   g93( wr_29   ,           wr_28   );
  nor   g94( wr_30   , wr_29   , wr_19   );
  not   g95( wr_31   ,           wr_30   );
  nor   g96( wr_32   , wr_31   , wr_17   );
  not   g97( wr_33   ,           wr_32   );
  nor   g98( wr_34   , wr_33   , wr_15   );
  not   g99( wr_35   ,           wr_34   );
  nor  g100( wr_36   , wr_35   , wr_13   );
  not  g101( wr_37   ,           wr_36   );
  nor  g102( wr_38   , wr_37   , wr_11   );
  not  g103( wr_39   ,           wr_38   );
  nor  g104( wr_41   , wr_38   , wr_9    );
  nor  g105( wr_40   , wr_39   , wr_9    );
  nor  g106( wr_44   , wr_43   , wr_41   );
  nor  g107( wr_117  , wr_116  , wr_41   );
  not  g108( G223gat ,           wr_40   );
  nor  g109( wr_59   , wr_40   , wr_58   );
  nor  g110( wr_66   , wr_40   , wr_65   );
  nor  g111( wr_73   , wr_40   , wr_72   );
  nor  g112( wr_80   , wr_40   , wr_79   );
  nor  g113( wr_87   , wr_40   , wr_86   );
  nor  g114( wr_94   , wr_40   , wr_93   );
  not  g115( wr_118  ,           wr_117  );
  nor  g116( wr_287  , wr_40   , wr_286  );
  nor  g117( wr_298  , wr_40   , wr_297  );
  nor  g118( wr_265  , wr_40   , wr_264  );
  nor  g119( wr_276  , wr_40   , wr_275  );
  nor  g120( wr_254  , wr_40   , wr_253  );
  nor  g121( wr_221  , wr_40   , wr_220  );
  nor  g122( wr_243  , wr_40   , wr_242  );
  nor  g123( wr_232  , wr_40   , wr_231  );
  nor  g124( wr_208  , wr_40   , wr_207  );
  nor  g125( wr_45   , G223gat , wr_11   );
  nor  g126( wr_51   , G223gat , wr_13   );
  nor  g127( wr_57   , G223gat , wr_15   );
  nor  g128( wr_64   , G223gat , wr_17   );
  nor  g129( wr_71   , G223gat , wr_19   );
  nor  g130( wr_78   , G223gat , wr_21   );
  nor  g131( wr_85   , G223gat , wr_23   );
  nor  g132( wr_92   , G223gat , wr_25   );
  nor  g133( wr_47   , wr_46   , wr_45   );
  nor  g134( wr_53   , wr_52   , wr_51   );
  nor  g135( wr_60   , wr_59   , wr_57   );
  nor  g136( wr_67   , wr_66   , wr_64   );
  nor  g137( wr_74   , wr_73   , wr_71   );
  nor  g138( wr_81   , wr_80   , wr_78   );
  nor  g139( wr_88   , wr_87   , wr_85   );
  nor  g140( wr_95   , wr_94   , wr_92   );
  nor  g141( wr_50   , wr_49   , wr_47   );
  nor  g142( wr_56   , wr_55   , wr_53   );
  nor  g143( wr_63   , wr_62   , wr_60   );
  nor  g144( wr_70   , wr_69   , wr_67   );
  nor  g145( wr_77   , wr_76   , wr_74   );
  nor  g146( wr_84   , wr_83   , wr_81   );
  nor  g147( wr_91   , wr_90   , wr_88   );
  nor  g148( wr_98   , wr_97   , wr_95   );
  nor  g149( wr_162  , wr_161  , wr_74   );
  nor  g150( wr_171  , wr_170  , wr_81   );
  nor  g151( wr_180  , wr_179  , wr_88   );
  nor  g152( wr_189  , wr_188  , wr_95   );
  nor  g153( wr_144  , wr_143  , wr_60   );
  nor  g154( wr_153  , wr_152  , wr_67   );
  nor  g155( wr_135  , wr_134  , wr_53   );
  nor  g156( wr_126  , wr_125  , wr_47   );
  nor  g157( wr_99   , wr_98   , wr_91   );
  not  g158( wr_139  ,           wr_63   );
  not  g159( wr_148  ,           wr_70   );
  not  g160( wr_154  ,           wr_153  );
  not  g161( wr_157  ,           wr_77   );
  not  g162( wr_163  ,           wr_162  );
  not  g163( wr_166  ,           wr_84   );
  not  g164( wr_172  ,           wr_171  );
  not  g165( wr_175  ,           wr_91   );
  not  g166( wr_181  ,           wr_180  );
  not  g167( wr_184  ,           wr_98   );
  not  g168( wr_190  ,           wr_189  );
  not  g169( wr_130  ,           wr_56   );
  not  g170( wr_145  ,           wr_144  );
  not  g171( wr_121  ,           wr_50   );
  not  g172( wr_136  ,           wr_135  );
  not  g173( wr_127  ,           wr_126  );
  not  g174( wr_100  ,           wr_99   );
  nor  g175( wr_101  , wr_100  , wr_84   );
  not  g176( wr_102  ,           wr_101  );
  nor  g177( wr_103  , wr_102  , wr_77   );
  not  g178( wr_104  ,           wr_103  );
  nor  g179( wr_105  , wr_104  , wr_70   );
  not  g180( wr_106  ,           wr_105  );
  nor  g181( wr_107  , wr_106  , wr_63   );
  not  g182( wr_108  ,           wr_107  );
  nor  g183( wr_109  , wr_108  , wr_56   );
  not  g184( wr_110  ,           wr_109  );
  nor  g185( wr_111  , wr_110  , wr_50   );
  not  g186( wr_112  ,           wr_111  );
  nor  g187( wr_114  , wr_111  , wr_44   );
  nor  g188( wr_113  , wr_112  , wr_44   );
  nor  g189( wr_119  , wr_118  , wr_114  );
  not  g190( G329gat ,           wr_113  );
  nor  g191( wr_158  , wr_113  , wr_157  );
  nor  g192( wr_167  , wr_113  , wr_166  );
  nor  g193( wr_176  , wr_113  , wr_175  );
  nor  g194( wr_185  , wr_113  , wr_184  );
  nor  g195( wr_140  , wr_113  , wr_139  );
  nor  g196( wr_149  , wr_113  , wr_148  );
  nor  g197( wr_131  , wr_113  , wr_130  );
  nor  g198( wr_122  , wr_113  , wr_121  );
  nor  g199( wr_285  , wr_113  , wr_284  );
  nor  g200( wr_296  , wr_113  , wr_295  );
  nor  g201( wr_263  , wr_113  , wr_262  );
  nor  g202( wr_274  , wr_113  , wr_273  );
  nor  g203( wr_252  , wr_113  , wr_251  );
  nor  g204( wr_219  , wr_113  , wr_218  );
  nor  g205( wr_241  , wr_113  , wr_240  );
  nor  g206( wr_212  , wr_113  , wr_211  );
  nor  g207( wr_230  , wr_113  , wr_229  );
  nor  g208( wr_156  , G329gat , wr_77   );
  nor  g209( wr_165  , G329gat , wr_84   );
  nor  g210( wr_174  , G329gat , wr_91   );
  nor  g211( wr_183  , G329gat , wr_98   );
  nor  g212( wr_138  , G329gat , wr_63   );
  nor  g213( wr_147  , G329gat , wr_70   );
  nor  g214( wr_129  , G329gat , wr_56   );
  nor  g215( wr_120  , G329gat , wr_50   );
  nor  g216( wr_150  , wr_149  , wr_147  );
  nor  g217( wr_159  , wr_158  , wr_156  );
  nor  g218( wr_168  , wr_167  , wr_165  );
  nor  g219( wr_177  , wr_176  , wr_174  );
  nor  g220( wr_186  , wr_185  , wr_183  );
  nor  g221( wr_141  , wr_140  , wr_138  );
  nor  g222( wr_132  , wr_131  , wr_129  );
  nor  g223( wr_123  , wr_122  , wr_120  );
  nor  g224( wr_173  , wr_172  , wr_168  );
  nor  g225( wr_182  , wr_181  , wr_177  );
  nor  g226( wr_191  , wr_190  , wr_186  );
  nor  g227( wr_155  , wr_154  , wr_150  );
  nor  g228( wr_164  , wr_163  , wr_159  );
  nor  g229( wr_146  , wr_145  , wr_141  );
  nor  g230( wr_137  , wr_136  , wr_132  );
  nor  g231( wr_128  , wr_127  , wr_123  );
  nor  g232( wr_192  , wr_191  , wr_182  );
  not  g233( wr_193  ,           wr_192  );
  nor  g234( wr_194  , wr_193  , wr_173  );
  not  g235( wr_195  ,           wr_194  );
  nor  g236( wr_196  , wr_195  , wr_164  );
  not  g237( wr_197  ,           wr_196  );
  nor  g238( wr_198  , wr_197  , wr_155  );
  not  g239( wr_199  ,           wr_198  );
  nor  g240( wr_200  , wr_199  , wr_146  );
  not  g241( wr_201  ,           wr_200  );
  nor  g242( wr_202  , wr_201  , wr_137  );
  not  g243( wr_203  ,           wr_202  );
  nor  g244( wr_204  , wr_203  , wr_128  );
  not  g245( wr_205  ,           wr_204  );
  nor  g246( wr_206  , wr_205  , wr_119  );
  nor  g247( wr_289  , wr_206  , wr_288  );
  nor  g248( wr_300  , wr_206  , wr_299  );
  nor  g249( wr_267  , wr_206  , wr_266  );
  nor  g250( wr_278  , wr_206  , wr_277  );
  nor  g251( wr_256  , wr_206  , wr_255  );
  nor  g252( wr_223  , wr_206  , wr_222  );
  nor  g253( wr_245  , wr_206  , wr_244  );
  nor  g254( wr_234  , wr_206  , wr_233  );
  nor  g255( wr_210  , wr_206  , wr_209  );
  not  g256( G370gat ,           wr_206  );
  nor  g257( wr_290  , wr_289  , wr_22   );
  nor  g258( wr_301  , wr_300  , wr_24   );
  nor  g259( wr_268  , wr_267  , wr_18   );
  nor  g260( wr_279  , wr_278  , wr_20   );
  nor  g261( wr_257  , wr_256  , wr_16   );
  nor  g262( wr_224  , wr_223  , wr_12   );
  nor  g263( wr_246  , wr_245  , wr_14   );
  nor  g264( wr_235  , wr_234  , wr_8    );
  nor  g265( wr_213  , wr_212  , wr_210  );
  not  g266( wr_291  ,           wr_290  );
  not  g267( wr_302  ,           wr_301  );
  not  g268( wr_269  ,           wr_268  );
  not  g269( wr_280  ,           wr_279  );
  not  g270( wr_258  ,           wr_257  );
  not  g271( wr_225  ,           wr_224  );
  not  g272( wr_247  ,           wr_246  );
  not  g273( wr_236  ,           wr_235  );
  not  g274( wr_214  ,           wr_213  );
  nor  g275( wr_292  , wr_291  , wr_287  );
  nor  g276( wr_303  , wr_302  , wr_298  );
  nor  g277( wr_270  , wr_269  , wr_265  );
  nor  g278( wr_281  , wr_280  , wr_276  );
  nor  g279( wr_259  , wr_258  , wr_254  );
  nor  g280( wr_226  , wr_225  , wr_221  );
  nor  g281( wr_248  , wr_247  , wr_243  );
  nor  g282( wr_237  , wr_236  , wr_232  );
  nor  g283( wr_215  , wr_214  , wr_10   );
  not  g284( wr_293  ,           wr_292  );
  not  g285( wr_304  ,           wr_303  );
  not  g286( wr_271  ,           wr_270  );
  not  g287( wr_282  ,           wr_281  );
  not  g288( wr_260  ,           wr_259  );
  not  g289( wr_227  ,           wr_226  );
  not  g290( wr_249  ,           wr_248  );
  not  g291( wr_238  ,           wr_237  );
  not  g292( wr_216  ,           wr_215  );
  nor  g293( wr_294  , wr_293  , wr_285  );
  nor  g294( wr_305  , wr_304  , wr_296  );
  nor  g295( wr_272  , wr_271  , wr_263  );
  nor  g296( wr_283  , wr_282  , wr_274  );
  nor  g297( wr_261  , wr_260  , wr_252  );
  nor  g298( wr_228  , wr_227  , wr_219  );
  nor  g299( wr_250  , wr_249  , wr_241  );
  nor  g300( wr_239  , wr_238  , wr_230  );
  nor  g301( wr_217  , wr_216  , wr_208  );
  nor  g302( wr_306  , wr_305  , wr_294  );
  not  g303( wr_330  ,           wr_272  );
  not  g304( wr_341  ,           wr_305  );
  not  g305( wr_326  ,           wr_283  );
  not  g306( wr_319  ,           wr_250  );
  not  g307( wr_307  ,           wr_306  );
  nor  g308( wr_331  , wr_330  , wr_261  );
  nor  g309( wr_342  , wr_341  , wr_283  );
  nor  g310( wr_327  , wr_326  , wr_261  );
  nor  g311( wr_320  , wr_319  , wr_228  );
  nor  g312( wr_308  , wr_307  , wr_283  );
  not  g313( wr_332  ,           wr_331  );
  not  g314( wr_343  ,           wr_342  );
  not  g315( wr_328  ,           wr_327  );
  nor  g316( wr_321  , wr_320  , wr_261  );
  not  g317( wr_309  ,           wr_308  );
  nor  g318( wr_333  , wr_332  , wr_228  );
  nor  g319( wr_344  , wr_343  , wr_228  );
  nor  g320( wr_329  , wr_328  , wr_250  );
  not  g321( wr_322  ,           wr_321  );
  nor  g322( wr_310  , wr_309  , wr_272  );
  not  g323( wr_334  ,           wr_333  );
  not  g324( wr_345  ,           wr_344  );
  nor  g325( wr_323  , wr_322  , wr_239  );
  not  g326( wr_311  ,           wr_310  );
  nor  g327( wr_335  , wr_334  , wr_250  );
  nor  g328( wr_346  , wr_345  , wr_250  );
  not  g329( wr_324  ,           wr_323  );
  nor  g330( wr_312  , wr_311  , wr_261  );
  nor  g331( wr_336  , wr_335  , wr_329  );
  nor  g332( wr_347  , wr_346  , wr_335  );
  nor  g333( wr_325  , wr_324  , wr_228  );
  not  g334( wr_313  ,           wr_312  );
  not  g335( wr_337  ,           wr_336  );
  not  g336( wr_348  ,           wr_347  );
  not  g337( G430gat ,           wr_325  );
  nor  g338( wr_314  , wr_313  , wr_250  );
  nor  g339( wr_338  , wr_337  , wr_239  );
  nor  g340( wr_349  , wr_348  , wr_239  );
  not  g341( wr_315  ,           wr_314  );
  not  g342( wr_339  ,           wr_338  );
  not  g343( wr_350  ,           wr_349  );
  nor  g344( wr_316  , wr_315  , wr_239  );
  nor  g345( wr_340  , wr_339  , wr_228  );
  nor  g346( wr_351  , wr_350  , wr_320  );
  not  g347( wr_317  ,           wr_316  );
  not  g348( G431gat ,           wr_340  );
  not  g349( G432gat ,           wr_351  );
  nor  g350( wr_318  , wr_317  , wr_228  );
  nor  g351( G421gat , wr_318  , wr_217  );

endmodule
