// Benchmark "./input/c1355" written by ABC on Thu Aug  8 02:45:58 2024

module c1355  ( 
    G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat,
    G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat,
    G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat,
    G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat,
    G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat,
    G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat,
    G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat,
    G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat,
    G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat,
    G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_G242gat_, new_G245gat_, new_G248gat_, new_G251gat_, new_G254gat_,
    new_G257gat_, new_G260gat_, new_G263gat_, new_G266gat_, new_G269gat_,
    new_G272gat_, new_G275gat_, new_G278gat_, new_G281gat_, new_G284gat_,
    new_G287gat_, new_G290gat_, new_G293gat_, new_G296gat_, new_G299gat_,
    new_G302gat_, new_G305gat_, new_G308gat_, new_G311gat_, new_G314gat_,
    new_G317gat_, new_G320gat_, new_G323gat_, new_G326gat_, new_G329gat_,
    new_G332gat_, new_G335gat_, new_G338gat_, new_G341gat_, new_G344gat_,
    new_G347gat_, new_G350gat_, new_G353gat_, new_G356gat_, new_G359gat_,
    new_G362gat_, new_G363gat_, new_G364gat_, new_G365gat_, new_G366gat_,
    new_G367gat_, new_G368gat_, new_G369gat_, new_G370gat_, new_G371gat_,
    new_G372gat_, new_G373gat_, new_G374gat_, new_G375gat_, new_G376gat_,
    new_G377gat_, new_G378gat_, new_G379gat_, new_G380gat_, new_G381gat_,
    new_G382gat_, new_G383gat_, new_G384gat_, new_G385gat_, new_G386gat_,
    new_G387gat_, new_G388gat_, new_G389gat_, new_G390gat_, new_G391gat_,
    new_G392gat_, new_G393gat_, new_G394gat_, new_G395gat_, new_G396gat_,
    new_G397gat_, new_G398gat_, new_G399gat_, new_G400gat_, new_G401gat_,
    new_G402gat_, new_G403gat_, new_G404gat_, new_G405gat_, new_G406gat_,
    new_G407gat_, new_G408gat_, new_G409gat_, new_G410gat_, new_G411gat_,
    new_G412gat_, new_G413gat_, new_G414gat_, new_G415gat_, new_G416gat_,
    new_G417gat_, new_G418gat_, new_G419gat_, new_G420gat_, new_G421gat_,
    new_G422gat_, new_G423gat_, new_G424gat_, new_G425gat_, new_G426gat_,
    new_G429gat_, new_G432gat_, new_G435gat_, new_G438gat_, new_G441gat_,
    new_G444gat_, new_G447gat_, new_G450gat_, new_G453gat_, new_G456gat_,
    new_G459gat_, new_G462gat_, new_G465gat_, new_G468gat_, new_G471gat_,
    new_G474gat_, new_G477gat_, new_G480gat_, new_G483gat_, new_G486gat_,
    new_G489gat_, new_G492gat_, new_G495gat_, new_G498gat_, new_G501gat_,
    new_G504gat_, new_G507gat_, new_G510gat_, new_G513gat_, new_G516gat_,
    new_G519gat_, new_G522gat_, new_G525gat_, new_G528gat_, new_G531gat_,
    new_G534gat_, new_G537gat_, new_G540gat_, new_G543gat_, new_G546gat_,
    new_G549gat_, new_G552gat_, new_G555gat_, new_G558gat_, new_G561gat_,
    new_G564gat_, new_G567gat_, new_G570gat_, new_G571gat_, new_G572gat_,
    new_G573gat_, new_G574gat_, new_G575gat_, new_G576gat_, new_G577gat_,
    new_G578gat_, new_G579gat_, new_G580gat_, new_G581gat_, new_G582gat_,
    new_G583gat_, new_G584gat_, new_G585gat_, new_G586gat_, new_G587gat_,
    new_G588gat_, new_G589gat_, new_G590gat_, new_G591gat_, new_G592gat_,
    new_G593gat_, new_G594gat_, new_G595gat_, new_G596gat_, new_G597gat_,
    new_G598gat_, new_G599gat_, new_G600gat_, new_G601gat_, new_G602gat_,
    new_G607gat_, new_G612gat_, new_G617gat_, new_G622gat_, new_G627gat_,
    new_G632gat_, new_G637gat_, new_G642gat_, new_G645gat_, new_G648gat_,
    new_G651gat_, new_G654gat_, new_G657gat_, new_G660gat_, new_G663gat_,
    new_G666gat_, new_G669gat_, new_G672gat_, new_G675gat_, new_G678gat_,
    new_G681gat_, new_G684gat_, new_G687gat_, new_G690gat_, new_G691gat_,
    new_G692gat_, new_G693gat_, new_G694gat_, new_G695gat_, new_G696gat_,
    new_G697gat_, new_G698gat_, new_G699gat_, new_G700gat_, new_G701gat_,
    new_G702gat_, new_G703gat_, new_G704gat_, new_G705gat_, new_G706gat_,
    new_G709gat_, new_G712gat_, new_G715gat_, new_G718gat_, new_G721gat_,
    new_G724gat_, new_G727gat_, new_G730gat_, new_G733gat_, new_G736gat_,
    new_G739gat_, new_G742gat_, new_G745gat_, new_G748gat_, new_G751gat_,
    new_G754gat_, new_G755gat_, new_G756gat_, new_G757gat_, new_G758gat_,
    new_G759gat_, new_G760gat_, new_G761gat_, new_G762gat_, new_G763gat_,
    new_G764gat_, new_G765gat_, new_G766gat_, new_G767gat_, new_G768gat_,
    new_G769gat_, new_G770gat_, new_G773gat_, new_G776gat_, new_G779gat_,
    new_G782gat_, new_G785gat_, new_G788gat_, new_G791gat_, new_G794gat_,
    new_G797gat_, new_G800gat_, new_G803gat_, new_G806gat_, new_G809gat_,
    new_G812gat_, new_G815gat_, new_G818gat_, new_G819gat_, new_G820gat_,
    new_G821gat_, new_G822gat_, new_G823gat_, new_G824gat_, new_G825gat_,
    new_G826gat_, new_G827gat_, new_G828gat_, new_G829gat_, new_G830gat_,
    new_G831gat_, new_G832gat_, new_G833gat_, new_G834gat_, new_G847gat_,
    new_G860gat_, new_G873gat_, new_G886gat_, new_G899gat_, new_G912gat_,
    new_G925gat_, new_G938gat_, new_G939gat_, new_G940gat_, new_G941gat_,
    new_G942gat_, new_G943gat_, new_G944gat_, new_G945gat_, new_G946gat_,
    new_G947gat_, new_G948gat_, new_G949gat_, new_G950gat_, new_G951gat_,
    new_G952gat_, new_G953gat_, new_G954gat_, new_G955gat_, new_G956gat_,
    new_G957gat_, new_G958gat_, new_G959gat_, new_G960gat_, new_G961gat_,
    new_G962gat_, new_G963gat_, new_G964gat_, new_G965gat_, new_G966gat_,
    new_G967gat_, new_G968gat_, new_G969gat_, new_G970gat_, new_G971gat_,
    new_G972gat_, new_G973gat_, new_G974gat_, new_G975gat_, new_G976gat_,
    new_G977gat_, new_G978gat_, new_G979gat_, new_G980gat_, new_G981gat_,
    new_G982gat_, new_G983gat_, new_G984gat_, new_G985gat_, new_G986gat_,
    new_G991gat_, new_G996gat_, new_G1001gat_, new_G1006gat_,
    new_G1011gat_, new_G1016gat_, new_G1021gat_, new_G1026gat_,
    new_G1031gat_, new_G1036gat_, new_G1039gat_, new_G1042gat_,
    new_G1045gat_, new_G1048gat_, new_G1051gat_, new_G1054gat_,
    new_G1057gat_, new_G1060gat_, new_G1063gat_, new_G1066gat_,
    new_G1069gat_, new_G1072gat_, new_G1075gat_, new_G1078gat_,
    new_G1081gat_, new_G1084gat_, new_G1087gat_, new_G1090gat_,
    new_G1093gat_, new_G1096gat_, new_G1099gat_, new_G1102gat_,
    new_G1105gat_, new_G1108gat_, new_G1111gat_, new_G1114gat_,
    new_G1117gat_, new_G1120gat_, new_G1123gat_, new_G1126gat_,
    new_G1129gat_, new_G1132gat_, new_G1135gat_, new_G1138gat_,
    new_G1141gat_, new_G1144gat_, new_G1147gat_, new_G1150gat_,
    new_G1153gat_, new_G1156gat_, new_G1159gat_, new_G1162gat_,
    new_G1165gat_, new_G1168gat_, new_G1171gat_, new_G1174gat_,
    new_G1177gat_, new_G1180gat_, new_G1183gat_, new_G1186gat_,
    new_G1189gat_, new_G1192gat_, new_G1195gat_, new_G1198gat_,
    new_G1201gat_, new_G1204gat_, new_G1207gat_, new_G1210gat_,
    new_G1213gat_, new_G1216gat_, new_G1219gat_, new_G1222gat_,
    new_G1225gat_, new_G1228gat_, new_G1229gat_, new_G1230gat_,
    new_G1231gat_, new_G1232gat_, new_G1233gat_, new_G1234gat_,
    new_G1235gat_, new_G1236gat_, new_G1237gat_, new_G1238gat_,
    new_G1239gat_, new_G1240gat_, new_G1241gat_, new_G1242gat_,
    new_G1243gat_, new_G1244gat_, new_G1245gat_, new_G1246gat_,
    new_G1247gat_, new_G1248gat_, new_G1249gat_, new_G1250gat_,
    new_G1251gat_, new_G1252gat_, new_G1253gat_, new_G1254gat_,
    new_G1255gat_, new_G1256gat_, new_G1257gat_, new_G1258gat_,
    new_G1259gat_, new_G1260gat_, new_G1261gat_, new_G1262gat_,
    new_G1263gat_, new_G1264gat_, new_G1265gat_, new_G1266gat_,
    new_G1267gat_, new_G1268gat_, new_G1269gat_, new_G1270gat_,
    new_G1271gat_, new_G1272gat_, new_G1273gat_, new_G1274gat_,
    new_G1275gat_, new_G1276gat_, new_G1277gat_, new_G1278gat_,
    new_G1279gat_, new_G1280gat_, new_G1281gat_, new_G1282gat_,
    new_G1283gat_, new_G1284gat_, new_G1285gat_, new_G1286gat_,
    new_G1287gat_, new_G1288gat_, new_G1289gat_, new_G1290gat_,
    new_G1291gat_, new_G1292gat_, new_G1293gat_, new_G1294gat_,
    new_G1295gat_, new_G1296gat_, new_G1297gat_, new_G1298gat_,
    new_G1299gat_, new_G1300gat_, new_G1301gat_, new_G1302gat_,
    new_G1303gat_, new_G1304gat_, new_G1305gat_, new_G1306gat_,
    new_G1307gat_, new_G1308gat_, new_G1309gat_, new_G1310gat_,
    new_G1311gat_, new_G1312gat_, new_G1313gat_, new_G1314gat_,
    new_G1315gat_, new_G1316gat_, new_G1317gat_, new_G1318gat_,
    new_G1319gat_, new_G1320gat_, new_G1321gat_, new_G1322gat_,
    new_G1323gat_;
  assign new_G242gat_ = G225gat & G233gat;
  assign new_G245gat_ = G226gat & G233gat;
  assign new_G248gat_ = G227gat & G233gat;
  assign new_G251gat_ = G228gat & G233gat;
  assign new_G254gat_ = G229gat & G233gat;
  assign new_G257gat_ = G230gat & G233gat;
  assign new_G260gat_ = G231gat & G233gat;
  assign new_G263gat_ = G232gat & G233gat;
  assign new_G266gat_ = ~G1gat | ~G8gat;
  assign new_G269gat_ = ~G15gat | ~G22gat;
  assign new_G272gat_ = ~G29gat | ~G36gat;
  assign new_G275gat_ = ~G43gat | ~G50gat;
  assign new_G278gat_ = ~G57gat | ~G64gat;
  assign new_G281gat_ = ~G71gat | ~G78gat;
  assign new_G284gat_ = ~G85gat | ~G92gat;
  assign new_G287gat_ = ~G99gat | ~G106gat;
  assign new_G290gat_ = ~G113gat | ~G120gat;
  assign new_G293gat_ = ~G127gat | ~G134gat;
  assign new_G296gat_ = ~G141gat | ~G148gat;
  assign new_G299gat_ = ~G155gat | ~G162gat;
  assign new_G302gat_ = ~G169gat | ~G176gat;
  assign new_G305gat_ = ~G183gat | ~G190gat;
  assign new_G308gat_ = ~G197gat | ~G204gat;
  assign new_G311gat_ = ~G211gat | ~G218gat;
  assign new_G314gat_ = ~G1gat | ~G29gat;
  assign new_G317gat_ = ~G57gat | ~G85gat;
  assign new_G320gat_ = ~G8gat | ~G36gat;
  assign new_G323gat_ = ~G64gat | ~G92gat;
  assign new_G326gat_ = ~G15gat | ~G43gat;
  assign new_G329gat_ = ~G71gat | ~G99gat;
  assign new_G332gat_ = ~G22gat | ~G50gat;
  assign new_G335gat_ = ~G78gat | ~G106gat;
  assign new_G338gat_ = ~G113gat | ~G141gat;
  assign new_G341gat_ = ~G169gat | ~G197gat;
  assign new_G344gat_ = ~G120gat | ~G148gat;
  assign new_G347gat_ = ~G176gat | ~G204gat;
  assign new_G350gat_ = ~G127gat | ~G155gat;
  assign new_G353gat_ = ~G183gat | ~G211gat;
  assign new_G356gat_ = ~G134gat | ~G162gat;
  assign new_G359gat_ = ~G190gat | ~G218gat;
  assign new_G362gat_ = ~G1gat | ~new_G266gat_;
  assign new_G363gat_ = ~G8gat | ~new_G266gat_;
  assign new_G364gat_ = ~G15gat | ~new_G269gat_;
  assign new_G365gat_ = ~G22gat | ~new_G269gat_;
  assign new_G366gat_ = ~G29gat | ~new_G272gat_;
  assign new_G367gat_ = ~G36gat | ~new_G272gat_;
  assign new_G368gat_ = ~G43gat | ~new_G275gat_;
  assign new_G369gat_ = ~G50gat | ~new_G275gat_;
  assign new_G370gat_ = ~G57gat | ~new_G278gat_;
  assign new_G371gat_ = ~G64gat | ~new_G278gat_;
  assign new_G372gat_ = ~G71gat | ~new_G281gat_;
  assign new_G373gat_ = ~G78gat | ~new_G281gat_;
  assign new_G374gat_ = ~G85gat | ~new_G284gat_;
  assign new_G375gat_ = ~G92gat | ~new_G284gat_;
  assign new_G376gat_ = ~G99gat | ~new_G287gat_;
  assign new_G377gat_ = ~G106gat | ~new_G287gat_;
  assign new_G378gat_ = ~G113gat | ~new_G290gat_;
  assign new_G379gat_ = ~G120gat | ~new_G290gat_;
  assign new_G380gat_ = ~G127gat | ~new_G293gat_;
  assign new_G381gat_ = ~G134gat | ~new_G293gat_;
  assign new_G382gat_ = ~G141gat | ~new_G296gat_;
  assign new_G383gat_ = ~G148gat | ~new_G296gat_;
  assign new_G384gat_ = ~G155gat | ~new_G299gat_;
  assign new_G385gat_ = ~G162gat | ~new_G299gat_;
  assign new_G386gat_ = ~G169gat | ~new_G302gat_;
  assign new_G387gat_ = ~G176gat | ~new_G302gat_;
  assign new_G388gat_ = ~G183gat | ~new_G305gat_;
  assign new_G389gat_ = ~G190gat | ~new_G305gat_;
  assign new_G390gat_ = ~G197gat | ~new_G308gat_;
  assign new_G391gat_ = ~G204gat | ~new_G308gat_;
  assign new_G392gat_ = ~G211gat | ~new_G311gat_;
  assign new_G393gat_ = ~G218gat | ~new_G311gat_;
  assign new_G394gat_ = ~G1gat | ~new_G314gat_;
  assign new_G395gat_ = ~G29gat | ~new_G314gat_;
  assign new_G396gat_ = ~G57gat | ~new_G317gat_;
  assign new_G397gat_ = ~G85gat | ~new_G317gat_;
  assign new_G398gat_ = ~G8gat | ~new_G320gat_;
  assign new_G399gat_ = ~G36gat | ~new_G320gat_;
  assign new_G400gat_ = ~G64gat | ~new_G323gat_;
  assign new_G401gat_ = ~G92gat | ~new_G323gat_;
  assign new_G402gat_ = ~G15gat | ~new_G326gat_;
  assign new_G403gat_ = ~G43gat | ~new_G326gat_;
  assign new_G404gat_ = ~G71gat | ~new_G329gat_;
  assign new_G405gat_ = ~G99gat | ~new_G329gat_;
  assign new_G406gat_ = ~G22gat | ~new_G332gat_;
  assign new_G407gat_ = ~G50gat | ~new_G332gat_;
  assign new_G408gat_ = ~G78gat | ~new_G335gat_;
  assign new_G409gat_ = ~G106gat | ~new_G335gat_;
  assign new_G410gat_ = ~G113gat | ~new_G338gat_;
  assign new_G411gat_ = ~G141gat | ~new_G338gat_;
  assign new_G412gat_ = ~G169gat | ~new_G341gat_;
  assign new_G413gat_ = ~G197gat | ~new_G341gat_;
  assign new_G414gat_ = ~G120gat | ~new_G344gat_;
  assign new_G415gat_ = ~G148gat | ~new_G344gat_;
  assign new_G416gat_ = ~G176gat | ~new_G347gat_;
  assign new_G417gat_ = ~G204gat | ~new_G347gat_;
  assign new_G418gat_ = ~G127gat | ~new_G350gat_;
  assign new_G419gat_ = ~G155gat | ~new_G350gat_;
  assign new_G420gat_ = ~G183gat | ~new_G353gat_;
  assign new_G421gat_ = ~G211gat | ~new_G353gat_;
  assign new_G422gat_ = ~G134gat | ~new_G356gat_;
  assign new_G423gat_ = ~G162gat | ~new_G356gat_;
  assign new_G424gat_ = ~G190gat | ~new_G359gat_;
  assign new_G425gat_ = ~G218gat | ~new_G359gat_;
  assign new_G426gat_ = ~new_G362gat_ | ~new_G363gat_;
  assign new_G429gat_ = ~new_G364gat_ | ~new_G365gat_;
  assign new_G432gat_ = ~new_G366gat_ | ~new_G367gat_;
  assign new_G435gat_ = ~new_G368gat_ | ~new_G369gat_;
  assign new_G438gat_ = ~new_G370gat_ | ~new_G371gat_;
  assign new_G441gat_ = ~new_G372gat_ | ~new_G373gat_;
  assign new_G444gat_ = ~new_G374gat_ | ~new_G375gat_;
  assign new_G447gat_ = ~new_G376gat_ | ~new_G377gat_;
  assign new_G450gat_ = ~new_G378gat_ | ~new_G379gat_;
  assign new_G453gat_ = ~new_G380gat_ | ~new_G381gat_;
  assign new_G456gat_ = ~new_G382gat_ | ~new_G383gat_;
  assign new_G459gat_ = ~new_G384gat_ | ~new_G385gat_;
  assign new_G462gat_ = ~new_G386gat_ | ~new_G387gat_;
  assign new_G465gat_ = ~new_G388gat_ | ~new_G389gat_;
  assign new_G468gat_ = ~new_G390gat_ | ~new_G391gat_;
  assign new_G471gat_ = ~new_G392gat_ | ~new_G393gat_;
  assign new_G474gat_ = ~new_G394gat_ | ~new_G395gat_;
  assign new_G477gat_ = ~new_G396gat_ | ~new_G397gat_;
  assign new_G480gat_ = ~new_G398gat_ | ~new_G399gat_;
  assign new_G483gat_ = ~new_G400gat_ | ~new_G401gat_;
  assign new_G486gat_ = ~new_G402gat_ | ~new_G403gat_;
  assign new_G489gat_ = ~new_G404gat_ | ~new_G405gat_;
  assign new_G492gat_ = ~new_G406gat_ | ~new_G407gat_;
  assign new_G495gat_ = ~new_G408gat_ | ~new_G409gat_;
  assign new_G498gat_ = ~new_G410gat_ | ~new_G411gat_;
  assign new_G501gat_ = ~new_G412gat_ | ~new_G413gat_;
  assign new_G504gat_ = ~new_G414gat_ | ~new_G415gat_;
  assign new_G507gat_ = ~new_G416gat_ | ~new_G417gat_;
  assign new_G510gat_ = ~new_G418gat_ | ~new_G419gat_;
  assign new_G513gat_ = ~new_G420gat_ | ~new_G421gat_;
  assign new_G516gat_ = ~new_G422gat_ | ~new_G423gat_;
  assign new_G519gat_ = ~new_G424gat_ | ~new_G425gat_;
  assign new_G522gat_ = ~new_G426gat_ | ~new_G429gat_;
  assign new_G525gat_ = ~new_G432gat_ | ~new_G435gat_;
  assign new_G528gat_ = ~new_G438gat_ | ~new_G441gat_;
  assign new_G531gat_ = ~new_G444gat_ | ~new_G447gat_;
  assign new_G534gat_ = ~new_G450gat_ | ~new_G453gat_;
  assign new_G537gat_ = ~new_G456gat_ | ~new_G459gat_;
  assign new_G540gat_ = ~new_G462gat_ | ~new_G465gat_;
  assign new_G543gat_ = ~new_G468gat_ | ~new_G471gat_;
  assign new_G546gat_ = ~new_G474gat_ | ~new_G477gat_;
  assign new_G549gat_ = ~new_G480gat_ | ~new_G483gat_;
  assign new_G552gat_ = ~new_G486gat_ | ~new_G489gat_;
  assign new_G555gat_ = ~new_G492gat_ | ~new_G495gat_;
  assign new_G558gat_ = ~new_G498gat_ | ~new_G501gat_;
  assign new_G561gat_ = ~new_G504gat_ | ~new_G507gat_;
  assign new_G564gat_ = ~new_G510gat_ | ~new_G513gat_;
  assign new_G567gat_ = ~new_G516gat_ | ~new_G519gat_;
  assign new_G570gat_ = ~new_G426gat_ | ~new_G522gat_;
  assign new_G571gat_ = ~new_G429gat_ | ~new_G522gat_;
  assign new_G572gat_ = ~new_G432gat_ | ~new_G525gat_;
  assign new_G573gat_ = ~new_G435gat_ | ~new_G525gat_;
  assign new_G574gat_ = ~new_G438gat_ | ~new_G528gat_;
  assign new_G575gat_ = ~new_G441gat_ | ~new_G528gat_;
  assign new_G576gat_ = ~new_G444gat_ | ~new_G531gat_;
  assign new_G577gat_ = ~new_G447gat_ | ~new_G531gat_;
  assign new_G578gat_ = ~new_G450gat_ | ~new_G534gat_;
  assign new_G579gat_ = ~new_G453gat_ | ~new_G534gat_;
  assign new_G580gat_ = ~new_G456gat_ | ~new_G537gat_;
  assign new_G581gat_ = ~new_G459gat_ | ~new_G537gat_;
  assign new_G582gat_ = ~new_G462gat_ | ~new_G540gat_;
  assign new_G583gat_ = ~new_G465gat_ | ~new_G540gat_;
  assign new_G584gat_ = ~new_G468gat_ | ~new_G543gat_;
  assign new_G585gat_ = ~new_G471gat_ | ~new_G543gat_;
  assign new_G586gat_ = ~new_G474gat_ | ~new_G546gat_;
  assign new_G587gat_ = ~new_G477gat_ | ~new_G546gat_;
  assign new_G588gat_ = ~new_G480gat_ | ~new_G549gat_;
  assign new_G589gat_ = ~new_G483gat_ | ~new_G549gat_;
  assign new_G590gat_ = ~new_G486gat_ | ~new_G552gat_;
  assign new_G591gat_ = ~new_G489gat_ | ~new_G552gat_;
  assign new_G592gat_ = ~new_G492gat_ | ~new_G555gat_;
  assign new_G593gat_ = ~new_G495gat_ | ~new_G555gat_;
  assign new_G594gat_ = ~new_G498gat_ | ~new_G558gat_;
  assign new_G595gat_ = ~new_G501gat_ | ~new_G558gat_;
  assign new_G596gat_ = ~new_G504gat_ | ~new_G561gat_;
  assign new_G597gat_ = ~new_G507gat_ | ~new_G561gat_;
  assign new_G598gat_ = ~new_G510gat_ | ~new_G564gat_;
  assign new_G599gat_ = ~new_G513gat_ | ~new_G564gat_;
  assign new_G600gat_ = ~new_G516gat_ | ~new_G567gat_;
  assign new_G601gat_ = ~new_G519gat_ | ~new_G567gat_;
  assign new_G602gat_ = ~new_G570gat_ | ~new_G571gat_;
  assign new_G607gat_ = ~new_G572gat_ | ~new_G573gat_;
  assign new_G612gat_ = ~new_G574gat_ | ~new_G575gat_;
  assign new_G617gat_ = ~new_G576gat_ | ~new_G577gat_;
  assign new_G622gat_ = ~new_G578gat_ | ~new_G579gat_;
  assign new_G627gat_ = ~new_G580gat_ | ~new_G581gat_;
  assign new_G632gat_ = ~new_G582gat_ | ~new_G583gat_;
  assign new_G637gat_ = ~new_G584gat_ | ~new_G585gat_;
  assign new_G642gat_ = ~new_G586gat_ | ~new_G587gat_;
  assign new_G645gat_ = ~new_G588gat_ | ~new_G589gat_;
  assign new_G648gat_ = ~new_G590gat_ | ~new_G591gat_;
  assign new_G651gat_ = ~new_G592gat_ | ~new_G593gat_;
  assign new_G654gat_ = ~new_G594gat_ | ~new_G595gat_;
  assign new_G657gat_ = ~new_G596gat_ | ~new_G597gat_;
  assign new_G660gat_ = ~new_G598gat_ | ~new_G599gat_;
  assign new_G663gat_ = ~new_G600gat_ | ~new_G601gat_;
  assign new_G666gat_ = ~new_G602gat_ | ~new_G607gat_;
  assign new_G669gat_ = ~new_G612gat_ | ~new_G617gat_;
  assign new_G672gat_ = ~new_G602gat_ | ~new_G612gat_;
  assign new_G675gat_ = ~new_G607gat_ | ~new_G617gat_;
  assign new_G678gat_ = ~new_G622gat_ | ~new_G627gat_;
  assign new_G681gat_ = ~new_G632gat_ | ~new_G637gat_;
  assign new_G684gat_ = ~new_G622gat_ | ~new_G632gat_;
  assign new_G687gat_ = ~new_G627gat_ | ~new_G637gat_;
  assign new_G690gat_ = ~new_G602gat_ | ~new_G666gat_;
  assign new_G691gat_ = ~new_G607gat_ | ~new_G666gat_;
  assign new_G692gat_ = ~new_G612gat_ | ~new_G669gat_;
  assign new_G693gat_ = ~new_G617gat_ | ~new_G669gat_;
  assign new_G694gat_ = ~new_G602gat_ | ~new_G672gat_;
  assign new_G695gat_ = ~new_G612gat_ | ~new_G672gat_;
  assign new_G696gat_ = ~new_G607gat_ | ~new_G675gat_;
  assign new_G697gat_ = ~new_G617gat_ | ~new_G675gat_;
  assign new_G698gat_ = ~new_G622gat_ | ~new_G678gat_;
  assign new_G699gat_ = ~new_G627gat_ | ~new_G678gat_;
  assign new_G700gat_ = ~new_G632gat_ | ~new_G681gat_;
  assign new_G701gat_ = ~new_G637gat_ | ~new_G681gat_;
  assign new_G702gat_ = ~new_G622gat_ | ~new_G684gat_;
  assign new_G703gat_ = ~new_G632gat_ | ~new_G684gat_;
  assign new_G704gat_ = ~new_G627gat_ | ~new_G687gat_;
  assign new_G705gat_ = ~new_G637gat_ | ~new_G687gat_;
  assign new_G706gat_ = ~new_G690gat_ | ~new_G691gat_;
  assign new_G709gat_ = ~new_G692gat_ | ~new_G693gat_;
  assign new_G712gat_ = ~new_G694gat_ | ~new_G695gat_;
  assign new_G715gat_ = ~new_G696gat_ | ~new_G697gat_;
  assign new_G718gat_ = ~new_G698gat_ | ~new_G699gat_;
  assign new_G721gat_ = ~new_G700gat_ | ~new_G701gat_;
  assign new_G724gat_ = ~new_G702gat_ | ~new_G703gat_;
  assign new_G727gat_ = ~new_G704gat_ | ~new_G705gat_;
  assign new_G730gat_ = ~new_G242gat_ | ~new_G718gat_;
  assign new_G733gat_ = ~new_G245gat_ | ~new_G721gat_;
  assign new_G736gat_ = ~new_G248gat_ | ~new_G724gat_;
  assign new_G739gat_ = ~new_G251gat_ | ~new_G727gat_;
  assign new_G742gat_ = ~new_G254gat_ | ~new_G706gat_;
  assign new_G745gat_ = ~new_G257gat_ | ~new_G709gat_;
  assign new_G748gat_ = ~new_G260gat_ | ~new_G712gat_;
  assign new_G751gat_ = ~new_G263gat_ | ~new_G715gat_;
  assign new_G754gat_ = ~new_G242gat_ | ~new_G730gat_;
  assign new_G755gat_ = ~new_G718gat_ | ~new_G730gat_;
  assign new_G756gat_ = ~new_G245gat_ | ~new_G733gat_;
  assign new_G757gat_ = ~new_G721gat_ | ~new_G733gat_;
  assign new_G758gat_ = ~new_G248gat_ | ~new_G736gat_;
  assign new_G759gat_ = ~new_G724gat_ | ~new_G736gat_;
  assign new_G760gat_ = ~new_G251gat_ | ~new_G739gat_;
  assign new_G761gat_ = ~new_G727gat_ | ~new_G739gat_;
  assign new_G762gat_ = ~new_G254gat_ | ~new_G742gat_;
  assign new_G763gat_ = ~new_G706gat_ | ~new_G742gat_;
  assign new_G764gat_ = ~new_G257gat_ | ~new_G745gat_;
  assign new_G765gat_ = ~new_G709gat_ | ~new_G745gat_;
  assign new_G766gat_ = ~new_G260gat_ | ~new_G748gat_;
  assign new_G767gat_ = ~new_G712gat_ | ~new_G748gat_;
  assign new_G768gat_ = ~new_G263gat_ | ~new_G751gat_;
  assign new_G769gat_ = ~new_G715gat_ | ~new_G751gat_;
  assign new_G770gat_ = ~new_G754gat_ | ~new_G755gat_;
  assign new_G773gat_ = ~new_G756gat_ | ~new_G757gat_;
  assign new_G776gat_ = ~new_G758gat_ | ~new_G759gat_;
  assign new_G779gat_ = ~new_G760gat_ | ~new_G761gat_;
  assign new_G782gat_ = ~new_G762gat_ | ~new_G763gat_;
  assign new_G785gat_ = ~new_G764gat_ | ~new_G765gat_;
  assign new_G788gat_ = ~new_G766gat_ | ~new_G767gat_;
  assign new_G791gat_ = ~new_G768gat_ | ~new_G769gat_;
  assign new_G794gat_ = ~new_G642gat_ | ~new_G770gat_;
  assign new_G797gat_ = ~new_G645gat_ | ~new_G773gat_;
  assign new_G800gat_ = ~new_G648gat_ | ~new_G776gat_;
  assign new_G803gat_ = ~new_G651gat_ | ~new_G779gat_;
  assign new_G806gat_ = ~new_G654gat_ | ~new_G782gat_;
  assign new_G809gat_ = ~new_G657gat_ | ~new_G785gat_;
  assign new_G812gat_ = ~new_G660gat_ | ~new_G788gat_;
  assign new_G815gat_ = ~new_G663gat_ | ~new_G791gat_;
  assign new_G818gat_ = ~new_G642gat_ | ~new_G794gat_;
  assign new_G819gat_ = ~new_G770gat_ | ~new_G794gat_;
  assign new_G820gat_ = ~new_G645gat_ | ~new_G797gat_;
  assign new_G821gat_ = ~new_G773gat_ | ~new_G797gat_;
  assign new_G822gat_ = ~new_G648gat_ | ~new_G800gat_;
  assign new_G823gat_ = ~new_G776gat_ | ~new_G800gat_;
  assign new_G824gat_ = ~new_G651gat_ | ~new_G803gat_;
  assign new_G825gat_ = ~new_G779gat_ | ~new_G803gat_;
  assign new_G826gat_ = ~new_G654gat_ | ~new_G806gat_;
  assign new_G827gat_ = ~new_G782gat_ | ~new_G806gat_;
  assign new_G828gat_ = ~new_G657gat_ | ~new_G809gat_;
  assign new_G829gat_ = ~new_G785gat_ | ~new_G809gat_;
  assign new_G830gat_ = ~new_G660gat_ | ~new_G812gat_;
  assign new_G831gat_ = ~new_G788gat_ | ~new_G812gat_;
  assign new_G832gat_ = ~new_G663gat_ | ~new_G815gat_;
  assign new_G833gat_ = ~new_G791gat_ | ~new_G815gat_;
  assign new_G834gat_ = ~new_G818gat_ | ~new_G819gat_;
  assign new_G847gat_ = ~new_G820gat_ | ~new_G821gat_;
  assign new_G860gat_ = ~new_G822gat_ | ~new_G823gat_;
  assign new_G873gat_ = ~new_G824gat_ | ~new_G825gat_;
  assign new_G886gat_ = ~new_G828gat_ | ~new_G829gat_;
  assign new_G899gat_ = ~new_G832gat_ | ~new_G833gat_;
  assign new_G912gat_ = ~new_G830gat_ | ~new_G831gat_;
  assign new_G925gat_ = ~new_G826gat_ | ~new_G827gat_;
  assign new_G938gat_ = ~new_G834gat_;
  assign new_G939gat_ = ~new_G847gat_;
  assign new_G940gat_ = ~new_G860gat_;
  assign new_G941gat_ = ~new_G834gat_;
  assign new_G942gat_ = ~new_G847gat_;
  assign new_G943gat_ = ~new_G873gat_;
  assign new_G944gat_ = ~new_G834gat_;
  assign new_G945gat_ = ~new_G860gat_;
  assign new_G946gat_ = ~new_G873gat_;
  assign new_G947gat_ = ~new_G847gat_;
  assign new_G948gat_ = ~new_G860gat_;
  assign new_G949gat_ = ~new_G873gat_;
  assign new_G950gat_ = ~new_G886gat_;
  assign new_G951gat_ = ~new_G899gat_;
  assign new_G952gat_ = ~new_G886gat_;
  assign new_G953gat_ = ~new_G912gat_;
  assign new_G954gat_ = ~new_G925gat_;
  assign new_G955gat_ = ~new_G899gat_;
  assign new_G956gat_ = ~new_G925gat_;
  assign new_G957gat_ = ~new_G912gat_;
  assign new_G958gat_ = ~new_G925gat_;
  assign new_G959gat_ = ~new_G886gat_;
  assign new_G960gat_ = ~new_G912gat_;
  assign new_G961gat_ = ~new_G925gat_;
  assign new_G962gat_ = ~new_G886gat_;
  assign new_G963gat_ = ~new_G899gat_;
  assign new_G964gat_ = ~new_G925gat_;
  assign new_G965gat_ = ~new_G912gat_;
  assign new_G966gat_ = ~new_G899gat_;
  assign new_G967gat_ = ~new_G886gat_;
  assign new_G968gat_ = ~new_G912gat_;
  assign new_G969gat_ = ~new_G899gat_;
  assign new_G970gat_ = ~new_G847gat_;
  assign new_G971gat_ = ~new_G873gat_;
  assign new_G972gat_ = ~new_G847gat_;
  assign new_G973gat_ = ~new_G860gat_;
  assign new_G974gat_ = ~new_G834gat_;
  assign new_G975gat_ = ~new_G873gat_;
  assign new_G976gat_ = ~new_G834gat_;
  assign new_G977gat_ = ~new_G860gat_;
  assign new_G978gat_ = new_G873gat_ & new_G940gat_ & new_G938gat_ & new_G939gat_;
  assign new_G979gat_ = new_G943gat_ & new_G860gat_ & new_G941gat_ & new_G942gat_;
  assign new_G980gat_ = new_G946gat_ & new_G945gat_ & new_G944gat_ & new_G847gat_;
  assign new_G981gat_ = new_G949gat_ & new_G948gat_ & new_G834gat_ & new_G947gat_;
  assign new_G982gat_ = new_G899gat_ & new_G960gat_ & new_G958gat_ & new_G959gat_;
  assign new_G983gat_ = new_G963gat_ & new_G912gat_ & new_G961gat_ & new_G962gat_;
  assign new_G984gat_ = new_G966gat_ & new_G965gat_ & new_G964gat_ & new_G886gat_;
  assign new_G985gat_ = new_G969gat_ & new_G968gat_ & new_G925gat_ & new_G967gat_;
  assign new_G986gat_ = new_G981gat_ | new_G980gat_ | new_G978gat_ | new_G979gat_;
  assign new_G991gat_ = new_G985gat_ | new_G984gat_ | new_G982gat_ | new_G983gat_;
  assign new_G996gat_ = new_G986gat_ & new_G951gat_ & new_G912gat_ & new_G925gat_ & new_G950gat_;
  assign new_G1001gat_ = new_G986gat_ & new_G899gat_ & new_G953gat_ & new_G925gat_ & new_G952gat_;
  assign new_G1006gat_ = new_G986gat_ & new_G955gat_ & new_G912gat_ & new_G954gat_ & new_G886gat_;
  assign new_G1011gat_ = new_G986gat_ & new_G899gat_ & new_G957gat_ & new_G956gat_ & new_G886gat_;
  assign new_G1016gat_ = new_G991gat_ & new_G971gat_ & new_G860gat_ & new_G834gat_ & new_G970gat_;
  assign new_G1021gat_ = new_G991gat_ & new_G873gat_ & new_G973gat_ & new_G834gat_ & new_G972gat_;
  assign new_G1026gat_ = new_G991gat_ & new_G975gat_ & new_G860gat_ & new_G974gat_ & new_G847gat_;
  assign new_G1031gat_ = new_G991gat_ & new_G873gat_ & new_G977gat_ & new_G976gat_ & new_G847gat_;
  assign new_G1036gat_ = new_G834gat_ & new_G996gat_;
  assign new_G1039gat_ = new_G847gat_ & new_G996gat_;
  assign new_G1042gat_ = new_G860gat_ & new_G996gat_;
  assign new_G1045gat_ = new_G873gat_ & new_G996gat_;
  assign new_G1048gat_ = new_G834gat_ & new_G1001gat_;
  assign new_G1051gat_ = new_G847gat_ & new_G1001gat_;
  assign new_G1054gat_ = new_G860gat_ & new_G1001gat_;
  assign new_G1057gat_ = new_G873gat_ & new_G1001gat_;
  assign new_G1060gat_ = new_G834gat_ & new_G1006gat_;
  assign new_G1063gat_ = new_G847gat_ & new_G1006gat_;
  assign new_G1066gat_ = new_G860gat_ & new_G1006gat_;
  assign new_G1069gat_ = new_G873gat_ & new_G1006gat_;
  assign new_G1072gat_ = new_G834gat_ & new_G1011gat_;
  assign new_G1075gat_ = new_G847gat_ & new_G1011gat_;
  assign new_G1078gat_ = new_G860gat_ & new_G1011gat_;
  assign new_G1081gat_ = new_G873gat_ & new_G1011gat_;
  assign new_G1084gat_ = new_G925gat_ & new_G1016gat_;
  assign new_G1087gat_ = new_G886gat_ & new_G1016gat_;
  assign new_G1090gat_ = new_G912gat_ & new_G1016gat_;
  assign new_G1093gat_ = new_G899gat_ & new_G1016gat_;
  assign new_G1096gat_ = new_G925gat_ & new_G1021gat_;
  assign new_G1099gat_ = new_G886gat_ & new_G1021gat_;
  assign new_G1102gat_ = new_G912gat_ & new_G1021gat_;
  assign new_G1105gat_ = new_G899gat_ & new_G1021gat_;
  assign new_G1108gat_ = new_G925gat_ & new_G1026gat_;
  assign new_G1111gat_ = new_G886gat_ & new_G1026gat_;
  assign new_G1114gat_ = new_G912gat_ & new_G1026gat_;
  assign new_G1117gat_ = new_G899gat_ & new_G1026gat_;
  assign new_G1120gat_ = new_G925gat_ & new_G1031gat_;
  assign new_G1123gat_ = new_G886gat_ & new_G1031gat_;
  assign new_G1126gat_ = new_G912gat_ & new_G1031gat_;
  assign new_G1129gat_ = new_G899gat_ & new_G1031gat_;
  assign new_G1132gat_ = ~G1gat | ~new_G1036gat_;
  assign new_G1135gat_ = ~G8gat | ~new_G1039gat_;
  assign new_G1138gat_ = ~G15gat | ~new_G1042gat_;
  assign new_G1141gat_ = ~G22gat | ~new_G1045gat_;
  assign new_G1144gat_ = ~G29gat | ~new_G1048gat_;
  assign new_G1147gat_ = ~G36gat | ~new_G1051gat_;
  assign new_G1150gat_ = ~G43gat | ~new_G1054gat_;
  assign new_G1153gat_ = ~G50gat | ~new_G1057gat_;
  assign new_G1156gat_ = ~G57gat | ~new_G1060gat_;
  assign new_G1159gat_ = ~G64gat | ~new_G1063gat_;
  assign new_G1162gat_ = ~G71gat | ~new_G1066gat_;
  assign new_G1165gat_ = ~G78gat | ~new_G1069gat_;
  assign new_G1168gat_ = ~G85gat | ~new_G1072gat_;
  assign new_G1171gat_ = ~G92gat | ~new_G1075gat_;
  assign new_G1174gat_ = ~G99gat | ~new_G1078gat_;
  assign new_G1177gat_ = ~G106gat | ~new_G1081gat_;
  assign new_G1180gat_ = ~G113gat | ~new_G1084gat_;
  assign new_G1183gat_ = ~G120gat | ~new_G1087gat_;
  assign new_G1186gat_ = ~G127gat | ~new_G1090gat_;
  assign new_G1189gat_ = ~G134gat | ~new_G1093gat_;
  assign new_G1192gat_ = ~G141gat | ~new_G1096gat_;
  assign new_G1195gat_ = ~G148gat | ~new_G1099gat_;
  assign new_G1198gat_ = ~G155gat | ~new_G1102gat_;
  assign new_G1201gat_ = ~G162gat | ~new_G1105gat_;
  assign new_G1204gat_ = ~G169gat | ~new_G1108gat_;
  assign new_G1207gat_ = ~G176gat | ~new_G1111gat_;
  assign new_G1210gat_ = ~G183gat | ~new_G1114gat_;
  assign new_G1213gat_ = ~G190gat | ~new_G1117gat_;
  assign new_G1216gat_ = ~G197gat | ~new_G1120gat_;
  assign new_G1219gat_ = ~G204gat | ~new_G1123gat_;
  assign new_G1222gat_ = ~G211gat | ~new_G1126gat_;
  assign new_G1225gat_ = ~G218gat | ~new_G1129gat_;
  assign new_G1228gat_ = ~G1gat | ~new_G1132gat_;
  assign new_G1229gat_ = ~new_G1036gat_ | ~new_G1132gat_;
  assign new_G1230gat_ = ~G8gat | ~new_G1135gat_;
  assign new_G1231gat_ = ~new_G1039gat_ | ~new_G1135gat_;
  assign new_G1232gat_ = ~G15gat | ~new_G1138gat_;
  assign new_G1233gat_ = ~new_G1042gat_ | ~new_G1138gat_;
  assign new_G1234gat_ = ~G22gat | ~new_G1141gat_;
  assign new_G1235gat_ = ~new_G1045gat_ | ~new_G1141gat_;
  assign new_G1236gat_ = ~G29gat | ~new_G1144gat_;
  assign new_G1237gat_ = ~new_G1048gat_ | ~new_G1144gat_;
  assign new_G1238gat_ = ~G36gat | ~new_G1147gat_;
  assign new_G1239gat_ = ~new_G1051gat_ | ~new_G1147gat_;
  assign new_G1240gat_ = ~G43gat | ~new_G1150gat_;
  assign new_G1241gat_ = ~new_G1054gat_ | ~new_G1150gat_;
  assign new_G1242gat_ = ~G50gat | ~new_G1153gat_;
  assign new_G1243gat_ = ~new_G1057gat_ | ~new_G1153gat_;
  assign new_G1244gat_ = ~G57gat | ~new_G1156gat_;
  assign new_G1245gat_ = ~new_G1060gat_ | ~new_G1156gat_;
  assign new_G1246gat_ = ~G64gat | ~new_G1159gat_;
  assign new_G1247gat_ = ~new_G1063gat_ | ~new_G1159gat_;
  assign new_G1248gat_ = ~G71gat | ~new_G1162gat_;
  assign new_G1249gat_ = ~new_G1066gat_ | ~new_G1162gat_;
  assign new_G1250gat_ = ~G78gat | ~new_G1165gat_;
  assign new_G1251gat_ = ~new_G1069gat_ | ~new_G1165gat_;
  assign new_G1252gat_ = ~G85gat | ~new_G1168gat_;
  assign new_G1253gat_ = ~new_G1072gat_ | ~new_G1168gat_;
  assign new_G1254gat_ = ~G92gat | ~new_G1171gat_;
  assign new_G1255gat_ = ~new_G1075gat_ | ~new_G1171gat_;
  assign new_G1256gat_ = ~G99gat | ~new_G1174gat_;
  assign new_G1257gat_ = ~new_G1078gat_ | ~new_G1174gat_;
  assign new_G1258gat_ = ~G106gat | ~new_G1177gat_;
  assign new_G1259gat_ = ~new_G1081gat_ | ~new_G1177gat_;
  assign new_G1260gat_ = ~G113gat | ~new_G1180gat_;
  assign new_G1261gat_ = ~new_G1084gat_ | ~new_G1180gat_;
  assign new_G1262gat_ = ~G120gat | ~new_G1183gat_;
  assign new_G1263gat_ = ~new_G1087gat_ | ~new_G1183gat_;
  assign new_G1264gat_ = ~G127gat | ~new_G1186gat_;
  assign new_G1265gat_ = ~new_G1090gat_ | ~new_G1186gat_;
  assign new_G1266gat_ = ~G134gat | ~new_G1189gat_;
  assign new_G1267gat_ = ~new_G1093gat_ | ~new_G1189gat_;
  assign new_G1268gat_ = ~G141gat | ~new_G1192gat_;
  assign new_G1269gat_ = ~new_G1096gat_ | ~new_G1192gat_;
  assign new_G1270gat_ = ~G148gat | ~new_G1195gat_;
  assign new_G1271gat_ = ~new_G1099gat_ | ~new_G1195gat_;
  assign new_G1272gat_ = ~G155gat | ~new_G1198gat_;
  assign new_G1273gat_ = ~new_G1102gat_ | ~new_G1198gat_;
  assign new_G1274gat_ = ~G162gat | ~new_G1201gat_;
  assign new_G1275gat_ = ~new_G1105gat_ | ~new_G1201gat_;
  assign new_G1276gat_ = ~G169gat | ~new_G1204gat_;
  assign new_G1277gat_ = ~new_G1108gat_ | ~new_G1204gat_;
  assign new_G1278gat_ = ~G176gat | ~new_G1207gat_;
  assign new_G1279gat_ = ~new_G1111gat_ | ~new_G1207gat_;
  assign new_G1280gat_ = ~G183gat | ~new_G1210gat_;
  assign new_G1281gat_ = ~new_G1114gat_ | ~new_G1210gat_;
  assign new_G1282gat_ = ~G190gat | ~new_G1213gat_;
  assign new_G1283gat_ = ~new_G1117gat_ | ~new_G1213gat_;
  assign new_G1284gat_ = ~G197gat | ~new_G1216gat_;
  assign new_G1285gat_ = ~new_G1120gat_ | ~new_G1216gat_;
  assign new_G1286gat_ = ~G204gat | ~new_G1219gat_;
  assign new_G1287gat_ = ~new_G1123gat_ | ~new_G1219gat_;
  assign new_G1288gat_ = ~G211gat | ~new_G1222gat_;
  assign new_G1289gat_ = ~new_G1126gat_ | ~new_G1222gat_;
  assign new_G1290gat_ = ~G218gat | ~new_G1225gat_;
  assign new_G1291gat_ = ~new_G1129gat_ | ~new_G1225gat_;
  assign new_G1292gat_ = ~new_G1228gat_ | ~new_G1229gat_;
  assign new_G1293gat_ = ~new_G1230gat_ | ~new_G1231gat_;
  assign new_G1294gat_ = ~new_G1232gat_ | ~new_G1233gat_;
  assign new_G1295gat_ = ~new_G1234gat_ | ~new_G1235gat_;
  assign new_G1296gat_ = ~new_G1236gat_ | ~new_G1237gat_;
  assign new_G1297gat_ = ~new_G1238gat_ | ~new_G1239gat_;
  assign new_G1298gat_ = ~new_G1240gat_ | ~new_G1241gat_;
  assign new_G1299gat_ = ~new_G1242gat_ | ~new_G1243gat_;
  assign new_G1300gat_ = ~new_G1244gat_ | ~new_G1245gat_;
  assign new_G1301gat_ = ~new_G1246gat_ | ~new_G1247gat_;
  assign new_G1302gat_ = ~new_G1248gat_ | ~new_G1249gat_;
  assign new_G1303gat_ = ~new_G1250gat_ | ~new_G1251gat_;
  assign new_G1304gat_ = ~new_G1252gat_ | ~new_G1253gat_;
  assign new_G1305gat_ = ~new_G1254gat_ | ~new_G1255gat_;
  assign new_G1306gat_ = ~new_G1256gat_ | ~new_G1257gat_;
  assign new_G1307gat_ = ~new_G1258gat_ | ~new_G1259gat_;
  assign new_G1308gat_ = ~new_G1260gat_ | ~new_G1261gat_;
  assign new_G1309gat_ = ~new_G1262gat_ | ~new_G1263gat_;
  assign new_G1310gat_ = ~new_G1264gat_ | ~new_G1265gat_;
  assign new_G1311gat_ = ~new_G1266gat_ | ~new_G1267gat_;
  assign new_G1312gat_ = ~new_G1268gat_ | ~new_G1269gat_;
  assign new_G1313gat_ = ~new_G1270gat_ | ~new_G1271gat_;
  assign new_G1314gat_ = ~new_G1272gat_ | ~new_G1273gat_;
  assign new_G1315gat_ = ~new_G1274gat_ | ~new_G1275gat_;
  assign new_G1316gat_ = ~new_G1276gat_ | ~new_G1277gat_;
  assign new_G1317gat_ = ~new_G1278gat_ | ~new_G1279gat_;
  assign new_G1318gat_ = ~new_G1280gat_ | ~new_G1281gat_;
  assign new_G1319gat_ = ~new_G1282gat_ | ~new_G1283gat_;
  assign new_G1320gat_ = ~new_G1284gat_ | ~new_G1285gat_;
  assign new_G1321gat_ = ~new_G1286gat_ | ~new_G1287gat_;
  assign new_G1322gat_ = ~new_G1288gat_ | ~new_G1289gat_;
  assign new_G1323gat_ = ~new_G1290gat_ | ~new_G1291gat_;
  assign G1324gat = new_G1292gat_;
  assign G1325gat = new_G1293gat_;
  assign G1326gat = new_G1294gat_;
  assign G1327gat = new_G1295gat_;
  assign G1328gat = new_G1296gat_;
  assign G1329gat = new_G1297gat_;
  assign G1330gat = new_G1298gat_;
  assign G1331gat = new_G1299gat_;
  assign G1332gat = new_G1300gat_;
  assign G1333gat = new_G1301gat_;
  assign G1334gat = new_G1302gat_;
  assign G1335gat = new_G1303gat_;
  assign G1336gat = new_G1304gat_;
  assign G1337gat = new_G1305gat_;
  assign G1338gat = new_G1306gat_;
  assign G1339gat = new_G1307gat_;
  assign G1340gat = new_G1308gat_;
  assign G1341gat = new_G1309gat_;
  assign G1342gat = new_G1310gat_;
  assign G1343gat = new_G1311gat_;
  assign G1344gat = new_G1312gat_;
  assign G1345gat = new_G1313gat_;
  assign G1346gat = new_G1314gat_;
  assign G1347gat = new_G1315gat_;
  assign G1348gat = new_G1316gat_;
  assign G1349gat = new_G1317gat_;
  assign G1350gat = new_G1318gat_;
  assign G1351gat = new_G1319gat_;
  assign G1352gat = new_G1320gat_;
  assign G1353gat = new_G1321gat_;
  assign G1354gat = new_G1322gat_;
  assign G1355gat = new_G1323gat_;
endmodule


