// Benchmark "./input/c1908" written by ABC on Thu Aug  8 02:45:58 2024

module c1908  ( 
    G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
    G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237,
    G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_G149_, new_G153_, new_G156_, new_G160_, new_G165_, new_G168_,
    new_G171_, new_G175_, new_G179_, new_G184_, new_G188_, new_G191_,
    new_G194_, new_G198_, new_G202_, new_G206_, new_G231_, new_G233_,
    new_G241_, new_G244_, new_G245_, new_G248_, new_G517_, new_G529_,
    new_G541_, new_G553_, new_G859_, new_G862_, new_G907_, new_G909_,
    new_G911_, new_G918_, new_G919_, new_G922_, new_G926_, new_G930_,
    new_G932_, new_G934_, new_G938_, new_G943_, new_G947_, new_G949_,
    new_G1506_, new_G1514_, new_G1522_, new_G1530_, new_G1538_, new_G1546_,
    new_G1554_, new_G1562_, new_G1570_, new_G1578_, new_G1586_, new_G1594_,
    new_G1602_, new_G1610_, new_G1618_, new_G1626_, new_G1512_, new_G1520_,
    new_G1528_, new_G1536_, new_G1544_, new_G1552_, new_G1560_, new_G1568_,
    new_G1576_, new_G1584_, new_G1592_, new_G1600_, new_G1608_, new_G1616_,
    new_G1624_, new_G1632_, new_G50_, new_G52_, new_G56_, new_G58_,
    new_G62_, new_G64_, new_G251_, new_G254_, new_G288_, new_G291_,
    new_G299_, new_G302_, new_G318_, new_G321_, new_G327_, new_G330_,
    new_G352_, new_G355_, new_G369_, new_G382_, new_G385_, new_G853_,
    new_G856_, new_G893_, new_G954_, new_G955_, new_G1050_, new_G1053_,
    new_G1176_, new_G1179_, new_G1197_, new_G1207_, new_G1222_, new_G1244_,
    new_G1278_, new_G1290_, new_G1300_, new_G1312_, new_G1332_, new_G1335_,
    new_G1442_, new_G1450_, new_G1458_, new_G1466_, new_G1474_, new_G1482_,
    new_G1490_, new_G1498_, new_G1634_, new_G1644_, new_G1657_, new_G1665_,
    new_G1697_, new_G1705_, new_G1713_, new_G1721_, new_G1745_, new_G1753_,
    new_G1785_, new_G1793_, new_G1814_, new_G1817_, new_G1830_, new_G1833_,
    new_G1841_, new_G1849_, new_G1854_, new_G1857_, new_G1870_, new_G1873_,
    new_G1878_, new_G1881_, new_G1642_, new_G1652_, new_G1056_, new_G1057_,
    new_G1182_, new_G1183_, new_G1211_, new_G1298_, new_G1320_, new_G1338_,
    new_G1339_, new_G457_, new_G459_, new_G482_, new_G487_, new_G492_,
    new_G505_, new_G1456_, new_G1448_, new_G1472_, new_G1464_, new_G1488_,
    new_G1480_, new_G1504_, new_G1496_, new_G956_, new_G967_, new_G978_,
    new_G979_, new_G980_, new_G1661_, new_G990_, new_G1669_, new_G1030_,
    new_G1701_, new_G1040_, new_G1709_, new_G1058_, new_G1717_, new_G1068_,
    new_G1725_, new_G1078_, new_G1090_, new_G1100_, new_G1749_, new_G1112_,
    new_G1757_, new_G1154_, new_G1789_, new_G1166_, new_G1797_, new_G1194_,
    new_G1201_, new_G1204_, new_G1820_, new_G1821_, new_G1230_, new_G1836_,
    new_G1837_, new_G1252_, new_G1256_, new_G1845_, new_G1268_, new_G1853_,
    new_G1860_, new_G1861_, new_G1286_, new_G1876_, new_G1877_, new_G1308_,
    new_G1884_, new_G1885_, new_G1654_, new_G1662_, new_G1694_, new_G1702_,
    new_G1710_, new_G1718_, new_G1726_, new_G1734_, new_G1742_, new_G1750_,
    new_G1782_, new_G1790_, new_G1838_, new_G1846_, new_G297_, new_G298_,
    new_G361_, new_G362_, new_G404_, new_G405_, new_G1225_, new_G1226_,
    new_G1247_, new_G1248_, new_G1281_, new_G1282_, new_G1303_, new_G1304_,
    new_G1315_, new_G1316_, new_G998_, new_G988_, new_G268_, new_G1038_,
    new_G1048_, new_G1076_, new_G1066_, new_G1098_, new_G1120_, new_G1174_,
    new_G363_, new_G1210_, new_G373_, new_G1276_, new_G406_, new_G565_,
    new_G566_, new_G614_, new_G615_, new_G958_, new_G969_, new_G1660_,
    new_G984_, new_G1668_, new_G994_, new_G1700_, new_G1034_, new_G1708_,
    new_G1044_, new_G1716_, new_G1062_, new_G1724_, new_G1072_, new_G1732_,
    new_G1086_, new_G1740_, new_G1748_, new_G1104_, new_G1108_, new_G1756_,
    new_G1116_, new_G1788_, new_G1158_, new_G1162_, new_G1796_, new_G1170_,
    new_G1200_, new_G1203_, new_G1227_, new_G1249_, new_G1844_, new_G1260_,
    new_G1264_, new_G1852_, new_G1272_, new_G1283_, new_G1305_, new_G1317_,
    new_G1410_, new_G1418_, new_G1426_, new_G1434_, new_G269_, new_G372_,
    new_G983_, new_G993_, new_G1033_, new_G1043_, new_G1061_, new_G1071_,
    new_G1103_, new_G1115_, new_G1157_, new_G1169_, new_G1184_, new_G1202_,
    new_G1259_, new_G1271_, new_G1322_, new_G374_, new_G396_, new_G1321_,
    new_G1424_, new_G1416_, new_G1440_, new_G1432_, new_G985_, new_G995_,
    new_G1035_, new_G1045_, new_G1063_, new_G1073_, new_G1105_, new_G1117_,
    new_G1159_, new_G1171_, new_G1212_, new_G1231_, new_G1232_, new_G1253_,
    new_G1254_, new_G1261_, new_G1273_, new_G1287_, new_G1288_, new_G1309_,
    new_G1310_, new_G1192_, new_G397_, new_G1330_, new_G1000_, new_G1010_,
    new_G1233_, new_G1255_, new_G1289_, new_G1311_, new_G1381_, new_G257_,
    new_G999_, new_G260_, new_G989_, new_G272_, new_G1039_, new_G294_,
    new_G1049_, new_G305_, new_G1077_, new_G308_, new_G1067_, new_G333_,
    new_G1121_, new_G358_, new_G1175_, new_G1220_, new_G388_, new_G1277_,
    new_G398_, new_G1109_, new_G1110_, new_G1163_, new_G1164_, new_G1234_,
    new_G1265_, new_G1266_, new_G1822_, new_G1862_, new_G1865_, new_G258_,
    new_G261_, new_G273_, new_G1018_, new_G1008_, new_G295_, new_G306_,
    new_G309_, new_G334_, new_G359_, new_G389_, new_G1385_, new_G1111_,
    new_G1165_, new_G1267_, new_G1886_, new_G259_, new_G262_, new_G274_,
    new_G296_, new_G307_, new_G310_, new_G335_, new_G360_, new_G1242_,
    new_G390_, new_G1828_, new_G1868_, new_G1869_, new_G1373_, new_G1798_,
    new_G1825_, new_G265_, new_G314_, new_G336_, new_G407_, new_G1293_,
    new_G1294_, new_G1892_, new_G1777_, new_G1889_, new_G410_, new_G1377_,
    new_G1804_, new_G1237_, new_G1829_, new_G1295_, new_G1670_, new_G1678_,
    new_G1729_, new_G1737_, new_G1761_, new_G1769_, new_G340_, new_G343_,
    new_G1781_, new_G1238_, new_G1325_, new_G1893_, new_G1340_, new_G1352_,
    new_G1673_, new_G1681_, new_G1801_, new_G1897_, new_G1905_, new_G391_,
    new_G1299_, new_G1676_, new_G1684_, new_G1081_, new_G1733_, new_G1093_,
    new_G1741_, new_G1765_, new_G1773_, new_G1239_, new_G1326_, new_G1894_,
    new_G1902_, new_G392_, new_G1360_, new_G1003_, new_G1677_, new_G1013_,
    new_G1685_, new_G1082_, new_G1094_, new_G1122_, new_G1134_, new_G1187_,
    new_G1805_, new_G1327_, new_G1901_, new_G1348_, new_G1909_, new_G1758_,
    new_G1766_, new_G377_, new_G1243_, new_G393_, new_G1004_, new_G1014_,
    new_G1083_, new_G1095_, new_G1188_, new_G1900_, new_G1344_, new_G1908_,
    new_G1356_, new_G1142_, new_G378_, new_G399_, new_G1331_, new_G1005_,
    new_G1015_, new_G1764_, new_G1126_, new_G1130_, new_G1772_, new_G1138_,
    new_G1189_, new_G1343_, new_G1355_, new_G324_, new_G1099_, new_G379_,
    new_G400_, new_G449_, new_G1087_, new_G1088_, new_G1125_, new_G1137_,
    new_G1345_, new_G1357_, new_G1397_, new_G277_, new_G1019_, new_G280_,
    new_G1009_, new_G325_, new_G364_, new_G1193_, new_G401_, new_G1089_,
    new_G1127_, new_G1139_, new_G278_, new_G281_, new_G326_, new_G365_,
    new_G413_, new_G1361_, new_G1401_, new_G445_, new_G1349_, new_G1350_,
    new_G1389_, new_G1493_, new_G1501_, new_G1689_, new_G279_, new_G282_,
    new_G346_, new_G1143_, new_G366_, new_G414_, new_G453_, new_G1131_,
    new_G1132_, new_G1351_, new_G1365_, new_G1405_, new_G285_, new_G347_,
    new_G367_, new_G415_, new_G1393_, new_G556_, new_G1505_, new_G559_,
    new_G1497_, new_G1693_, new_G1133_, new_G1477_, new_G1485_, new_G1809_,
    new_G348_, new_G1369_, new_G1409_, new_G557_, new_G560_, new_G1362_,
    new_G1378_, new_G1429_, new_G1437_, new_G1686_, new_G1774_, new_G1910_,
    new_G1918_, new_G544_, new_G1489_, new_G547_, new_G1481_, new_G558_,
    new_G561_, new_G1813_, new_G1370_, new_G1368_, new_G417_, new_G1384_,
    new_G424_, new_G508_, new_G1441_, new_G511_, new_G1433_, new_G545_,
    new_G548_, new_G564_, new_G1692_, new_G1024_, new_G1780_, new_G1148_,
    new_G1916_, new_G1924_, new_G416_, new_G1376_, new_G421_, new_G423_,
    new_G509_, new_G512_, new_G546_, new_G549_, new_G719_, new_G722_,
    new_G1023_, new_G1147_, new_G418_, new_G420_, new_G425_, new_G510_,
    new_G513_, new_G552_, new_G1025_, new_G1149_, new_G419_, new_G422_,
    new_G441_, new_G516_, new_G725_, new_G728_, new_G1029_, new_G1153_,
    new_G433_, new_G437_, new_G663_, new_G666_, new_G731_, new_G746_,
    new_G756_, new_G770_, new_G1461_, new_G1469_, new_G1413_, new_G1421_,
    new_G1445_, new_G1453_, new_G532_, new_G1473_, new_G535_, new_G1465_,
    new_G495_, new_G1425_, new_G498_, new_G1417_, new_G520_, new_G1457_,
    new_G523_, new_G1449_, new_G533_, new_G536_, new_G496_, new_G499_,
    new_G521_, new_G524_, new_G534_, new_G537_, new_G497_, new_G500_,
    new_G522_, new_G525_, new_G540_, new_G503_, new_G528_, new_G669_,
    new_G672_, new_G569_, new_G588_, new_G618_, new_G639_, new_G867_,
    new_G588a_, new_G588b_, new_G639a_, new_G639b_, new_G675_, new_G688_,
    new_G696_, new_G710_, new_G73_, new_G572_, new_G573_, new_G621_,
    new_G622_, new_G776_, new_G780_, new_G784_, new_G788_, new_G812_,
    new_G832_, new_G836_, new_G1509_, new_G1517_, new_G1525_, new_G1533_,
    new_G1581_, new_G1621_, new_G1629_, new_G792_, new_G796_, new_G800_,
    new_G804_, new_G808_, new_G816_, new_G820_, new_G824_, new_G828_,
    new_G871_, new_G873_, new_G875_, new_G877_, new_G879_, new_G881_,
    new_G883_, new_G885_, new_G1541_, new_G1549_, new_G1557_, new_G1565_,
    new_G1573_, new_G1589_, new_G1597_, new_G1605_, new_G1613_, new_G1_,
    new_G1513_, new_G4_, new_G1521_, new_G7_, new_G1529_, new_G10_,
    new_G1537_, new_G28_, new_G1585_, new_G43_, new_G1625_, new_G46_,
    new_G1633_, new_G886_, new_G2_, new_G5_, new_G8_, new_G11_, new_G13_,
    new_G1545_, new_G16_, new_G1553_, new_G19_, new_G1561_, new_G22_,
    new_G1569_, new_G25_, new_G1577_, new_G29_, new_G31_, new_G1593_,
    new_G34_, new_G1601_, new_G37_, new_G1609_, new_G40_, new_G1617_,
    new_G44_, new_G47_, new_G857_, new_G860_, new_G863_, new_G865_,
    new_G14_, new_G17_, new_G20_, new_G23_, new_G26_, new_G32_, new_G35_,
    new_G38_, new_G41_, new_G1913_, new_G1921_, new_G887_, new_G462_,
    new_G74_, new_G1637_, new_G1917_, new_G1647_, new_G1925_, new_G1020_,
    new_G1144_, new_G1386_, new_G1394_, new_G1402_, new_G1638_, new_G1648_,
    new_G1806_, new_G1639_, new_G1649_, new_G287_, new_G350_, new_G427_,
    new_G429_, new_G431_, new_G1028_, new_G1152_, new_G1392_, new_G1400_,
    new_G1408_, new_G1812_, new_G1216_, new_G286_, new_G349_, new_G426_,
    new_G428_, new_G430_, new_G67_, new_G1643_, new_G70_, new_G1653_,
    new_G1215_, new_G49_, new_G53_, new_G59_, new_G61_, new_G65_, new_G68_,
    new_G71_, new_G1217_, new_G375_, new_G1221_, new_G376_, new_G55_;
  assign new_G149_ = ~G101;
  assign new_G153_ = ~G104;
  assign new_G156_ = ~G107;
  assign new_G160_ = ~G110;
  assign new_G165_ = ~G113;
  assign new_G168_ = ~G116;
  assign new_G171_ = ~G119;
  assign new_G175_ = ~G122;
  assign new_G179_ = ~G125;
  assign new_G184_ = ~G128;
  assign new_G188_ = ~G131;
  assign new_G191_ = ~G134;
  assign new_G194_ = ~G137;
  assign new_G198_ = ~G140;
  assign new_G202_ = ~G143;
  assign new_G206_ = ~G146;
  assign new_G231_ = ~G224 | ~G898;
  assign new_G233_ = ~G227 | ~G900;
  assign new_G241_ = ~G237;
  assign new_G244_ = ~G237;
  assign new_G245_ = G234;
  assign new_G248_ = G234;
  assign new_G517_ = ~G469;
  assign new_G529_ = ~G472;
  assign new_G541_ = ~G475;
  assign new_G553_ = ~G478;
  assign new_G859_ = ~G953;
  assign new_G862_ = ~G953;
  assign new_G907_ = ~G898;
  assign new_G909_ = ~G900;
  assign new_G911_ = G902;
  assign new_G918_ = ~G902;
  assign new_G919_ = G902;
  assign new_G922_ = ~G902;
  assign new_G926_ = G952;
  assign new_G930_ = ~G952;
  assign new_G932_ = ~G952;
  assign new_G934_ = G953;
  assign new_G938_ = ~G953;
  assign new_G943_ = G953;
  assign new_G947_ = G953;
  assign new_G949_ = ~G953;
  assign new_G1506_ = G101;
  assign new_G1514_ = G104;
  assign new_G1522_ = G107;
  assign new_G1530_ = G110;
  assign new_G1538_ = G113;
  assign new_G1546_ = G116;
  assign new_G1554_ = G119;
  assign new_G1562_ = G122;
  assign new_G1570_ = G125;
  assign new_G1578_ = G128;
  assign new_G1586_ = G131;
  assign new_G1594_ = G134;
  assign new_G1602_ = G137;
  assign new_G1610_ = G140;
  assign new_G1618_ = G143;
  assign new_G1626_ = G146;
  assign new_G1512_ = ~new_G1506_;
  assign new_G1520_ = ~new_G1514_;
  assign new_G1528_ = ~new_G1522_;
  assign new_G1536_ = ~new_G1530_;
  assign new_G1544_ = ~new_G1538_;
  assign new_G1552_ = ~new_G1546_;
  assign new_G1560_ = ~new_G1554_;
  assign new_G1568_ = ~new_G1562_;
  assign new_G1576_ = ~new_G1570_;
  assign new_G1584_ = ~new_G1578_;
  assign new_G1592_ = ~new_G1586_;
  assign new_G1600_ = ~new_G1594_;
  assign new_G1608_ = ~new_G1602_;
  assign new_G1616_ = ~new_G1610_;
  assign new_G1624_ = ~new_G1618_;
  assign new_G1632_ = ~new_G1626_;
  assign new_G50_ = ~new_G930_ | ~new_G947_;
  assign new_G52_ = ~new_G930_ | ~new_G947_;
  assign new_G56_ = ~new_G930_ | ~new_G947_;
  assign new_G58_ = ~new_G930_ | ~new_G947_;
  assign new_G62_ = ~new_G930_ | ~new_G947_;
  assign new_G64_ = ~new_G930_ | ~new_G947_;
  assign new_G251_ = new_G149_;
  assign new_G254_ = new_G153_;
  assign new_G288_ = new_G165_;
  assign new_G291_ = new_G168_;
  assign new_G299_ = new_G184_;
  assign new_G302_ = new_G202_;
  assign new_G318_ = G224 & new_G938_;
  assign new_G321_ = new_G179_;
  assign new_G327_ = new_G188_;
  assign new_G330_ = new_G191_;
  assign new_G352_ = G227 & new_G938_;
  assign new_G355_ = new_G198_;
  assign new_G369_ = new_G938_ & G210 & new_G241_;
  assign new_G382_ = new_G206_;
  assign new_G385_ = new_G198_;
  assign new_G853_ = ~new_G943_ | ~new_G907_;
  assign new_G856_ = ~new_G943_ | ~new_G909_;
  assign new_G893_ = ~new_G248_ | ~G237;
  assign new_G954_ = ~new_G248_ | ~new_G922_;
  assign new_G955_ = ~new_G244_ | ~new_G922_;
  assign new_G1050_ = new_G160_;
  assign new_G1053_ = new_G175_;
  assign new_G1176_ = new_G179_;
  assign new_G1179_ = new_G198_;
  assign new_G1197_ = new_G149_;
  assign new_G1207_ = new_G149_;
  assign new_G1222_ = new_G153_;
  assign new_G1244_ = new_G188_;
  assign new_G1278_ = new_G156_;
  assign new_G1290_ = new_G938_ & G217 & new_G245_;
  assign new_G1300_ = new_G191_;
  assign new_G1312_ = new_G160_;
  assign new_G1332_ = new_G194_;
  assign new_G1335_ = new_G938_ & G221 & new_G245_;
  assign new_G1442_ = new_G517_;
  assign new_G1450_ = new_G517_;
  assign new_G1458_ = new_G529_;
  assign new_G1466_ = new_G529_;
  assign new_G1474_ = new_G541_;
  assign new_G1482_ = new_G541_;
  assign new_G1490_ = new_G553_;
  assign new_G1498_ = new_G553_;
  assign new_G1634_ = new_G231_ & new_G934_;
  assign new_G1644_ = new_G233_ & new_G934_;
  assign new_G1657_ = new_G156_;
  assign new_G1665_ = new_G156_;
  assign new_G1697_ = new_G171_;
  assign new_G1705_ = new_G171_;
  assign new_G1713_ = new_G206_;
  assign new_G1721_ = new_G206_;
  assign new_G1745_ = new_G194_;
  assign new_G1753_ = new_G194_;
  assign new_G1785_ = new_G160_;
  assign new_G1793_ = new_G160_;
  assign new_G1814_ = new_G165_;
  assign new_G1817_ = new_G175_;
  assign new_G1830_ = new_G938_ & G214 & new_G241_;
  assign new_G1833_ = new_G202_;
  assign new_G1841_ = new_G179_;
  assign new_G1849_ = new_G179_;
  assign new_G1854_ = new_G168_;
  assign new_G1857_ = new_G175_;
  assign new_G1870_ = new_G184_;
  assign new_G1873_ = new_G202_;
  assign new_G1878_ = new_G171_;
  assign new_G1881_ = new_G184_;
  assign new_G1642_ = ~new_G1634_;
  assign new_G1652_ = ~new_G1644_;
  assign new_G1056_ = ~new_G1050_;
  assign new_G1057_ = ~new_G1053_;
  assign new_G1182_ = ~new_G1176_;
  assign new_G1183_ = ~new_G1179_;
  assign new_G1211_ = ~new_G1207_;
  assign new_G1298_ = ~new_G1290_;
  assign new_G1320_ = ~new_G1312_;
  assign new_G1338_ = ~new_G1332_;
  assign new_G1339_ = ~new_G1335_;
  assign new_G457_ = G210 & new_G955_;
  assign new_G459_ = G217 & new_G954_;
  assign new_G482_ = ~G214 | ~new_G955_;
  assign new_G487_ = ~G221 | ~new_G954_;
  assign new_G492_ = ~G210 | ~new_G955_;
  assign new_G505_ = ~G217 | ~new_G954_;
  assign new_G1456_ = ~new_G1450_;
  assign new_G1448_ = ~new_G1442_;
  assign new_G1472_ = ~new_G1466_;
  assign new_G1464_ = ~new_G1458_;
  assign new_G1488_ = ~new_G1482_;
  assign new_G1480_ = ~new_G1474_;
  assign new_G1504_ = ~new_G1498_;
  assign new_G1496_ = ~new_G1490_;
  assign new_G956_ = ~new_G893_ | ~new_G943_ | ~new_G907_ | ~new_G919_;
  assign new_G967_ = ~new_G893_ | ~new_G943_ | ~new_G909_ | ~new_G919_;
  assign new_G978_ = ~new_G893_ | ~new_G926_ | ~new_G949_;
  assign new_G979_ = new_G893_ & new_G926_ & new_G949_;
  assign new_G980_ = new_G251_;
  assign new_G1661_ = ~new_G1657_;
  assign new_G990_ = new_G251_;
  assign new_G1669_ = ~new_G1665_;
  assign new_G1030_ = new_G288_;
  assign new_G1701_ = ~new_G1697_;
  assign new_G1040_ = new_G288_;
  assign new_G1709_ = ~new_G1705_;
  assign new_G1058_ = new_G299_;
  assign new_G1717_ = ~new_G1713_;
  assign new_G1068_ = new_G299_;
  assign new_G1725_ = ~new_G1721_;
  assign new_G1078_ = new_G318_;
  assign new_G1090_ = new_G318_;
  assign new_G1100_ = new_G327_;
  assign new_G1749_ = ~new_G1745_;
  assign new_G1112_ = new_G327_;
  assign new_G1757_ = ~new_G1753_;
  assign new_G1154_ = new_G352_;
  assign new_G1789_ = ~new_G1785_;
  assign new_G1166_ = new_G352_;
  assign new_G1797_ = ~new_G1793_;
  assign new_G1194_ = new_G369_;
  assign new_G1201_ = ~new_G1197_;
  assign new_G1204_ = new_G369_;
  assign new_G1820_ = ~new_G1814_;
  assign new_G1821_ = ~new_G1817_;
  assign new_G1230_ = ~new_G1222_;
  assign new_G1836_ = ~new_G1830_;
  assign new_G1837_ = ~new_G1833_;
  assign new_G1252_ = ~new_G1244_;
  assign new_G1256_ = new_G382_;
  assign new_G1845_ = ~new_G1841_;
  assign new_G1268_ = new_G382_;
  assign new_G1853_ = ~new_G1849_;
  assign new_G1860_ = ~new_G1854_;
  assign new_G1861_ = ~new_G1857_;
  assign new_G1286_ = ~new_G1278_;
  assign new_G1876_ = ~new_G1870_;
  assign new_G1877_ = ~new_G1873_;
  assign new_G1308_ = ~new_G1300_;
  assign new_G1884_ = ~new_G1878_;
  assign new_G1885_ = ~new_G1881_;
  assign new_G1654_ = new_G254_;
  assign new_G1662_ = new_G254_;
  assign new_G1694_ = new_G291_;
  assign new_G1702_ = new_G291_;
  assign new_G1710_ = new_G302_;
  assign new_G1718_ = new_G302_;
  assign new_G1726_ = new_G321_;
  assign new_G1734_ = new_G321_;
  assign new_G1742_ = new_G330_;
  assign new_G1750_ = new_G330_;
  assign new_G1782_ = new_G355_;
  assign new_G1790_ = new_G355_;
  assign new_G1838_ = new_G385_;
  assign new_G1846_ = new_G385_;
  assign new_G297_ = ~new_G1053_ | ~new_G1056_;
  assign new_G298_ = ~new_G1050_ | ~new_G1057_;
  assign new_G361_ = ~new_G1179_ | ~new_G1182_;
  assign new_G362_ = ~new_G1176_ | ~new_G1183_;
  assign new_G404_ = ~new_G1335_ | ~new_G1338_;
  assign new_G405_ = ~new_G1332_ | ~new_G1339_;
  assign new_G1225_ = ~new_G1817_ | ~new_G1820_;
  assign new_G1226_ = ~new_G1814_ | ~new_G1821_;
  assign new_G1247_ = ~new_G1833_ | ~new_G1836_;
  assign new_G1248_ = ~new_G1830_ | ~new_G1837_;
  assign new_G1281_ = ~new_G1857_ | ~new_G1860_;
  assign new_G1282_ = ~new_G1854_ | ~new_G1861_;
  assign new_G1303_ = ~new_G1873_ | ~new_G1876_;
  assign new_G1304_ = ~new_G1870_ | ~new_G1877_;
  assign new_G1315_ = ~new_G1881_ | ~new_G1884_;
  assign new_G1316_ = ~new_G1878_ | ~new_G1885_;
  assign new_G998_ = ~new_G990_;
  assign new_G988_ = ~new_G980_;
  assign new_G268_ = ~new_G297_ | ~new_G298_;
  assign new_G1038_ = ~new_G1030_;
  assign new_G1048_ = ~new_G1040_;
  assign new_G1076_ = ~new_G1068_;
  assign new_G1066_ = ~new_G1058_;
  assign new_G1098_ = ~new_G1090_;
  assign new_G1120_ = ~new_G1112_;
  assign new_G1174_ = ~new_G1166_;
  assign new_G363_ = ~new_G361_ | ~new_G362_;
  assign new_G1210_ = ~new_G1204_;
  assign new_G373_ = ~new_G1204_ | ~new_G1211_;
  assign new_G1276_ = ~new_G1268_;
  assign new_G406_ = ~new_G404_ | ~new_G405_;
  assign new_G565_ = ~new_G482_;
  assign new_G566_ = new_G482_;
  assign new_G614_ = ~new_G487_;
  assign new_G615_ = new_G487_;
  assign new_G958_ = ~new_G956_ | ~new_G978_;
  assign new_G969_ = ~new_G967_ | ~new_G978_;
  assign new_G1660_ = ~new_G1654_;
  assign new_G984_ = ~new_G1654_ | ~new_G1661_;
  assign new_G1668_ = ~new_G1662_;
  assign new_G994_ = ~new_G1662_ | ~new_G1669_;
  assign new_G1700_ = ~new_G1694_;
  assign new_G1034_ = ~new_G1694_ | ~new_G1701_;
  assign new_G1708_ = ~new_G1702_;
  assign new_G1044_ = ~new_G1702_ | ~new_G1709_;
  assign new_G1716_ = ~new_G1710_;
  assign new_G1062_ = ~new_G1710_ | ~new_G1717_;
  assign new_G1724_ = ~new_G1718_;
  assign new_G1072_ = ~new_G1718_ | ~new_G1725_;
  assign new_G1732_ = ~new_G1726_;
  assign new_G1086_ = ~new_G1078_;
  assign new_G1740_ = ~new_G1734_;
  assign new_G1748_ = ~new_G1742_;
  assign new_G1104_ = ~new_G1742_ | ~new_G1749_;
  assign new_G1108_ = ~new_G1100_;
  assign new_G1756_ = ~new_G1750_;
  assign new_G1116_ = ~new_G1750_ | ~new_G1757_;
  assign new_G1788_ = ~new_G1782_;
  assign new_G1158_ = ~new_G1782_ | ~new_G1789_;
  assign new_G1162_ = ~new_G1154_;
  assign new_G1796_ = ~new_G1790_;
  assign new_G1170_ = ~new_G1790_ | ~new_G1797_;
  assign new_G1200_ = ~new_G1194_;
  assign new_G1203_ = ~new_G1194_ | ~new_G1201_;
  assign new_G1227_ = ~new_G1225_ | ~new_G1226_;
  assign new_G1249_ = ~new_G1247_ | ~new_G1248_;
  assign new_G1844_ = ~new_G1838_;
  assign new_G1260_ = ~new_G1838_ | ~new_G1845_;
  assign new_G1264_ = ~new_G1256_;
  assign new_G1852_ = ~new_G1846_;
  assign new_G1272_ = ~new_G1846_ | ~new_G1853_;
  assign new_G1283_ = ~new_G1281_ | ~new_G1282_;
  assign new_G1305_ = ~new_G1303_ | ~new_G1304_;
  assign new_G1317_ = ~new_G1315_ | ~new_G1316_;
  assign new_G1410_ = new_G492_;
  assign new_G1418_ = new_G492_;
  assign new_G1426_ = new_G505_;
  assign new_G1434_ = new_G505_;
  assign new_G269_ = ~new_G268_;
  assign new_G372_ = ~new_G1207_ | ~new_G1210_;
  assign new_G983_ = ~new_G1657_ | ~new_G1660_;
  assign new_G993_ = ~new_G1665_ | ~new_G1668_;
  assign new_G1033_ = ~new_G1697_ | ~new_G1700_;
  assign new_G1043_ = ~new_G1705_ | ~new_G1708_;
  assign new_G1061_ = ~new_G1713_ | ~new_G1716_;
  assign new_G1071_ = ~new_G1721_ | ~new_G1724_;
  assign new_G1103_ = ~new_G1745_ | ~new_G1748_;
  assign new_G1115_ = ~new_G1753_ | ~new_G1756_;
  assign new_G1157_ = ~new_G1785_ | ~new_G1788_;
  assign new_G1169_ = ~new_G1793_ | ~new_G1796_;
  assign new_G1184_ = ~new_G363_;
  assign new_G1202_ = ~new_G1197_ | ~new_G1200_;
  assign new_G1259_ = ~new_G1841_ | ~new_G1844_;
  assign new_G1271_ = ~new_G1849_ | ~new_G1852_;
  assign new_G1322_ = ~new_G406_;
  assign new_G374_ = ~new_G372_ | ~new_G373_;
  assign new_G396_ = ~new_G1317_ | ~new_G1320_;
  assign new_G1321_ = ~new_G1317_;
  assign new_G1424_ = ~new_G1418_;
  assign new_G1416_ = ~new_G1410_;
  assign new_G1440_ = ~new_G1434_;
  assign new_G1432_ = ~new_G1426_;
  assign new_G985_ = ~new_G983_ | ~new_G984_;
  assign new_G995_ = ~new_G993_ | ~new_G994_;
  assign new_G1035_ = ~new_G1033_ | ~new_G1034_;
  assign new_G1045_ = ~new_G1043_ | ~new_G1044_;
  assign new_G1063_ = ~new_G1061_ | ~new_G1062_;
  assign new_G1073_ = ~new_G1071_ | ~new_G1072_;
  assign new_G1105_ = ~new_G1103_ | ~new_G1104_;
  assign new_G1117_ = ~new_G1115_ | ~new_G1116_;
  assign new_G1159_ = ~new_G1157_ | ~new_G1158_;
  assign new_G1171_ = ~new_G1169_ | ~new_G1170_;
  assign new_G1212_ = ~new_G1202_ | ~new_G1203_;
  assign new_G1231_ = ~new_G1227_;
  assign new_G1232_ = ~new_G1227_ | ~new_G1230_;
  assign new_G1253_ = ~new_G1249_;
  assign new_G1254_ = ~new_G1249_ | ~new_G1252_;
  assign new_G1261_ = ~new_G1259_ | ~new_G1260_;
  assign new_G1273_ = ~new_G1271_ | ~new_G1272_;
  assign new_G1287_ = ~new_G1283_;
  assign new_G1288_ = ~new_G1283_ | ~new_G1286_;
  assign new_G1309_ = ~new_G1305_;
  assign new_G1310_ = ~new_G1305_ | ~new_G1308_;
  assign new_G1192_ = ~new_G1184_;
  assign new_G397_ = ~new_G1312_ | ~new_G1321_;
  assign new_G1330_ = ~new_G1322_;
  assign new_G1000_ = new_G269_;
  assign new_G1010_ = new_G269_;
  assign new_G1233_ = ~new_G1222_ | ~new_G1231_;
  assign new_G1255_ = ~new_G1244_ | ~new_G1253_;
  assign new_G1289_ = ~new_G1278_ | ~new_G1287_;
  assign new_G1311_ = ~new_G1300_ | ~new_G1309_;
  assign new_G1381_ = ~new_G374_;
  assign new_G257_ = ~new_G995_ | ~new_G998_;
  assign new_G999_ = ~new_G995_;
  assign new_G260_ = ~new_G985_ | ~new_G988_;
  assign new_G989_ = ~new_G985_;
  assign new_G272_ = ~new_G1035_ | ~new_G1038_;
  assign new_G1039_ = ~new_G1035_;
  assign new_G294_ = ~new_G1045_ | ~new_G1048_;
  assign new_G1049_ = ~new_G1045_;
  assign new_G305_ = ~new_G1073_ | ~new_G1076_;
  assign new_G1077_ = ~new_G1073_;
  assign new_G308_ = ~new_G1063_ | ~new_G1066_;
  assign new_G1067_ = ~new_G1063_;
  assign new_G333_ = ~new_G1117_ | ~new_G1120_;
  assign new_G1121_ = ~new_G1117_;
  assign new_G358_ = ~new_G1171_ | ~new_G1174_;
  assign new_G1175_ = ~new_G1171_;
  assign new_G1220_ = ~new_G1212_;
  assign new_G388_ = ~new_G1273_ | ~new_G1276_;
  assign new_G1277_ = ~new_G1273_;
  assign new_G398_ = ~new_G396_ | ~new_G397_;
  assign new_G1109_ = ~new_G1105_;
  assign new_G1110_ = ~new_G1105_ | ~new_G1108_;
  assign new_G1163_ = ~new_G1159_;
  assign new_G1164_ = ~new_G1159_ | ~new_G1162_;
  assign new_G1234_ = ~new_G1232_ | ~new_G1233_;
  assign new_G1265_ = ~new_G1261_;
  assign new_G1266_ = ~new_G1261_ | ~new_G1264_;
  assign new_G1822_ = ~new_G1254_ | ~new_G1255_;
  assign new_G1862_ = ~new_G1310_ | ~new_G1311_;
  assign new_G1865_ = ~new_G1288_ | ~new_G1289_;
  assign new_G258_ = ~new_G990_ | ~new_G999_;
  assign new_G261_ = ~new_G980_ | ~new_G989_;
  assign new_G273_ = ~new_G1030_ | ~new_G1039_;
  assign new_G1018_ = ~new_G1010_;
  assign new_G1008_ = ~new_G1000_;
  assign new_G295_ = ~new_G1040_ | ~new_G1049_;
  assign new_G306_ = ~new_G1068_ | ~new_G1077_;
  assign new_G309_ = ~new_G1058_ | ~new_G1067_;
  assign new_G334_ = ~new_G1112_ | ~new_G1121_;
  assign new_G359_ = ~new_G1166_ | ~new_G1175_;
  assign new_G389_ = ~new_G1268_ | ~new_G1277_;
  assign new_G1385_ = ~new_G1381_;
  assign new_G1111_ = ~new_G1100_ | ~new_G1109_;
  assign new_G1165_ = ~new_G1154_ | ~new_G1163_;
  assign new_G1267_ = ~new_G1256_ | ~new_G1265_;
  assign new_G1886_ = ~new_G398_;
  assign new_G259_ = ~new_G257_ | ~new_G258_;
  assign new_G262_ = ~new_G260_ | ~new_G261_;
  assign new_G274_ = ~new_G272_ | ~new_G273_;
  assign new_G296_ = ~new_G294_ | ~new_G295_;
  assign new_G307_ = ~new_G305_ | ~new_G306_;
  assign new_G310_ = ~new_G308_ | ~new_G309_;
  assign new_G335_ = ~new_G333_ | ~new_G334_;
  assign new_G360_ = ~new_G358_ | ~new_G359_;
  assign new_G1242_ = ~new_G1234_;
  assign new_G390_ = ~new_G388_ | ~new_G389_;
  assign new_G1828_ = ~new_G1822_;
  assign new_G1868_ = ~new_G1862_;
  assign new_G1869_ = ~new_G1865_;
  assign new_G1373_ = ~new_G1164_ | ~new_G1165_;
  assign new_G1798_ = ~new_G1110_ | ~new_G1111_;
  assign new_G1825_ = ~new_G1266_ | ~new_G1267_;
  assign new_G265_ = ~new_G259_;
  assign new_G314_ = ~new_G307_;
  assign new_G336_ = ~new_G335_;
  assign new_G407_ = ~new_G296_;
  assign new_G1293_ = ~new_G1865_ | ~new_G1868_;
  assign new_G1294_ = ~new_G1862_ | ~new_G1869_;
  assign new_G1892_ = ~new_G1886_;
  assign new_G1777_ = ~new_G360_;
  assign new_G1889_ = ~new_G390_;
  assign new_G410_ = new_G310_;
  assign new_G1377_ = ~new_G1373_;
  assign new_G1804_ = ~new_G1798_;
  assign new_G1237_ = ~new_G1825_ | ~new_G1828_;
  assign new_G1829_ = ~new_G1825_;
  assign new_G1295_ = ~new_G1293_ | ~new_G1294_;
  assign new_G1670_ = new_G274_;
  assign new_G1678_ = new_G274_;
  assign new_G1729_ = new_G310_;
  assign new_G1737_ = new_G310_;
  assign new_G1761_ = new_G262_;
  assign new_G1769_ = new_G262_;
  assign new_G340_ = new_G336_;
  assign new_G343_ = new_G314_;
  assign new_G1781_ = ~new_G1777_;
  assign new_G1238_ = ~new_G1822_ | ~new_G1829_;
  assign new_G1325_ = ~new_G1889_ | ~new_G1892_;
  assign new_G1893_ = ~new_G1889_;
  assign new_G1340_ = new_G407_;
  assign new_G1352_ = new_G407_;
  assign new_G1673_ = new_G265_;
  assign new_G1681_ = new_G265_;
  assign new_G1801_ = new_G314_;
  assign new_G1897_ = new_G336_;
  assign new_G1905_ = new_G336_;
  assign new_G391_ = ~new_G1295_ | ~new_G1298_;
  assign new_G1299_ = ~new_G1295_;
  assign new_G1676_ = ~new_G1670_;
  assign new_G1684_ = ~new_G1678_;
  assign new_G1081_ = ~new_G1729_ | ~new_G1732_;
  assign new_G1733_ = ~new_G1729_;
  assign new_G1093_ = ~new_G1737_ | ~new_G1740_;
  assign new_G1741_ = ~new_G1737_;
  assign new_G1765_ = ~new_G1761_;
  assign new_G1773_ = ~new_G1769_;
  assign new_G1239_ = ~new_G1237_ | ~new_G1238_;
  assign new_G1326_ = ~new_G1886_ | ~new_G1893_;
  assign new_G1894_ = new_G410_;
  assign new_G1902_ = new_G410_;
  assign new_G392_ = ~new_G1290_ | ~new_G1299_;
  assign new_G1360_ = ~new_G1352_;
  assign new_G1003_ = ~new_G1673_ | ~new_G1676_;
  assign new_G1677_ = ~new_G1673_;
  assign new_G1013_ = ~new_G1681_ | ~new_G1684_;
  assign new_G1685_ = ~new_G1681_;
  assign new_G1082_ = ~new_G1726_ | ~new_G1733_;
  assign new_G1094_ = ~new_G1734_ | ~new_G1741_;
  assign new_G1122_ = new_G340_;
  assign new_G1134_ = new_G340_;
  assign new_G1187_ = ~new_G1801_ | ~new_G1804_;
  assign new_G1805_ = ~new_G1801_;
  assign new_G1327_ = ~new_G1325_ | ~new_G1326_;
  assign new_G1901_ = ~new_G1897_;
  assign new_G1348_ = ~new_G1340_;
  assign new_G1909_ = ~new_G1905_;
  assign new_G1758_ = new_G343_;
  assign new_G1766_ = new_G343_;
  assign new_G377_ = ~new_G1239_ | ~new_G1242_;
  assign new_G1243_ = ~new_G1239_;
  assign new_G393_ = ~new_G391_ | ~new_G392_;
  assign new_G1004_ = ~new_G1670_ | ~new_G1677_;
  assign new_G1014_ = ~new_G1678_ | ~new_G1685_;
  assign new_G1083_ = ~new_G1081_ | ~new_G1082_;
  assign new_G1095_ = ~new_G1093_ | ~new_G1094_;
  assign new_G1188_ = ~new_G1798_ | ~new_G1805_;
  assign new_G1900_ = ~new_G1894_;
  assign new_G1344_ = ~new_G1894_ | ~new_G1901_;
  assign new_G1908_ = ~new_G1902_;
  assign new_G1356_ = ~new_G1902_ | ~new_G1909_;
  assign new_G1142_ = ~new_G1134_;
  assign new_G378_ = ~new_G1234_ | ~new_G1243_;
  assign new_G399_ = ~new_G1327_ | ~new_G1330_;
  assign new_G1331_ = ~new_G1327_;
  assign new_G1005_ = ~new_G1003_ | ~new_G1004_;
  assign new_G1015_ = ~new_G1013_ | ~new_G1014_;
  assign new_G1764_ = ~new_G1758_;
  assign new_G1126_ = ~new_G1758_ | ~new_G1765_;
  assign new_G1130_ = ~new_G1122_;
  assign new_G1772_ = ~new_G1766_;
  assign new_G1138_ = ~new_G1766_ | ~new_G1773_;
  assign new_G1189_ = ~new_G1187_ | ~new_G1188_;
  assign new_G1343_ = ~new_G1897_ | ~new_G1900_;
  assign new_G1355_ = ~new_G1905_ | ~new_G1908_;
  assign new_G324_ = ~new_G1095_ | ~new_G1098_;
  assign new_G1099_ = ~new_G1095_;
  assign new_G379_ = ~new_G377_ | ~new_G378_;
  assign new_G400_ = ~new_G1322_ | ~new_G1331_;
  assign new_G449_ = ~new_G393_ | ~new_G918_;
  assign new_G1087_ = ~new_G1083_;
  assign new_G1088_ = ~new_G1083_ | ~new_G1086_;
  assign new_G1125_ = ~new_G1761_ | ~new_G1764_;
  assign new_G1137_ = ~new_G1769_ | ~new_G1772_;
  assign new_G1345_ = ~new_G1343_ | ~new_G1344_;
  assign new_G1357_ = ~new_G1355_ | ~new_G1356_;
  assign new_G1397_ = new_G393_;
  assign new_G277_ = ~new_G1015_ | ~new_G1018_;
  assign new_G1019_ = ~new_G1015_;
  assign new_G280_ = ~new_G1005_ | ~new_G1008_;
  assign new_G1009_ = ~new_G1005_;
  assign new_G325_ = ~new_G1090_ | ~new_G1099_;
  assign new_G364_ = ~new_G1189_ | ~new_G1192_;
  assign new_G1193_ = ~new_G1189_;
  assign new_G401_ = ~new_G399_ | ~new_G400_;
  assign new_G1089_ = ~new_G1078_ | ~new_G1087_;
  assign new_G1127_ = ~new_G1125_ | ~new_G1126_;
  assign new_G1139_ = ~new_G1137_ | ~new_G1138_;
  assign new_G278_ = ~new_G1010_ | ~new_G1019_;
  assign new_G281_ = ~new_G1000_ | ~new_G1009_;
  assign new_G326_ = ~new_G324_ | ~new_G325_;
  assign new_G365_ = ~new_G1184_ | ~new_G1193_;
  assign new_G413_ = ~new_G1357_ | ~new_G1360_;
  assign new_G1361_ = ~new_G1357_;
  assign new_G1401_ = ~new_G1397_;
  assign new_G445_ = ~new_G379_ | ~new_G918_;
  assign new_G1349_ = ~new_G1345_;
  assign new_G1350_ = ~new_G1345_ | ~new_G1348_;
  assign new_G1389_ = new_G379_;
  assign new_G1493_ = new_G449_;
  assign new_G1501_ = new_G449_;
  assign new_G1689_ = ~new_G1088_ | ~new_G1089_;
  assign new_G279_ = ~new_G277_ | ~new_G278_;
  assign new_G282_ = ~new_G280_ | ~new_G281_;
  assign new_G346_ = ~new_G1139_ | ~new_G1142_;
  assign new_G1143_ = ~new_G1139_;
  assign new_G366_ = ~new_G364_ | ~new_G365_;
  assign new_G414_ = ~new_G1352_ | ~new_G1361_;
  assign new_G453_ = ~new_G401_ | ~new_G918_;
  assign new_G1131_ = ~new_G1127_;
  assign new_G1132_ = ~new_G1127_ | ~new_G1130_;
  assign new_G1351_ = ~new_G1340_ | ~new_G1349_;
  assign new_G1365_ = ~new_G326_;
  assign new_G1405_ = new_G401_;
  assign new_G285_ = ~new_G279_;
  assign new_G347_ = ~new_G1134_ | ~new_G1143_;
  assign new_G367_ = ~new_G366_;
  assign new_G415_ = ~new_G413_ | ~new_G414_;
  assign new_G1393_ = ~new_G1389_;
  assign new_G556_ = ~new_G1501_ | ~new_G1504_;
  assign new_G1505_ = ~new_G1501_;
  assign new_G559_ = ~new_G1493_ | ~new_G1496_;
  assign new_G1497_ = ~new_G1493_;
  assign new_G1693_ = ~new_G1689_;
  assign new_G1133_ = ~new_G1122_ | ~new_G1131_;
  assign new_G1477_ = new_G445_;
  assign new_G1485_ = new_G445_;
  assign new_G1809_ = ~new_G1350_ | ~new_G1351_;
  assign new_G348_ = ~new_G346_ | ~new_G347_;
  assign new_G1369_ = ~new_G1365_;
  assign new_G1409_ = ~new_G1405_;
  assign new_G557_ = ~new_G1498_ | ~new_G1505_;
  assign new_G560_ = ~new_G1490_ | ~new_G1497_;
  assign new_G1362_ = new_G282_;
  assign new_G1378_ = ~new_G415_;
  assign new_G1429_ = new_G453_;
  assign new_G1437_ = new_G453_;
  assign new_G1686_ = new_G282_;
  assign new_G1774_ = ~new_G1132_ | ~new_G1133_;
  assign new_G1910_ = new_G285_ & new_G853_;
  assign new_G1918_ = new_G856_ & new_G367_;
  assign new_G544_ = ~new_G1485_ | ~new_G1488_;
  assign new_G1489_ = ~new_G1485_;
  assign new_G547_ = ~new_G1477_ | ~new_G1480_;
  assign new_G1481_ = ~new_G1477_;
  assign new_G558_ = ~new_G556_ | ~new_G557_;
  assign new_G561_ = ~new_G559_ | ~new_G560_;
  assign new_G1813_ = ~new_G1809_;
  assign new_G1370_ = ~new_G348_;
  assign new_G1368_ = ~new_G1362_;
  assign new_G417_ = ~new_G1362_ | ~new_G1369_;
  assign new_G1384_ = ~new_G1378_;
  assign new_G424_ = ~new_G1378_ | ~new_G1385_;
  assign new_G508_ = ~new_G1437_ | ~new_G1440_;
  assign new_G1441_ = ~new_G1437_;
  assign new_G511_ = ~new_G1429_ | ~new_G1432_;
  assign new_G1433_ = ~new_G1429_;
  assign new_G545_ = ~new_G1482_ | ~new_G1489_;
  assign new_G548_ = ~new_G1474_ | ~new_G1481_;
  assign new_G564_ = ~new_G558_;
  assign new_G1692_ = ~new_G1686_;
  assign new_G1024_ = ~new_G1686_ | ~new_G1693_;
  assign new_G1780_ = ~new_G1774_;
  assign new_G1148_ = ~new_G1774_ | ~new_G1781_;
  assign new_G1916_ = ~new_G1910_;
  assign new_G1924_ = ~new_G1918_;
  assign new_G416_ = ~new_G1365_ | ~new_G1368_;
  assign new_G1376_ = ~new_G1370_;
  assign new_G421_ = ~new_G1370_ | ~new_G1377_;
  assign new_G423_ = ~new_G1381_ | ~new_G1384_;
  assign new_G509_ = ~new_G1434_ | ~new_G1441_;
  assign new_G512_ = ~new_G1426_ | ~new_G1433_;
  assign new_G546_ = ~new_G544_ | ~new_G545_;
  assign new_G549_ = ~new_G547_ | ~new_G548_;
  assign new_G719_ = ~new_G561_;
  assign new_G722_ = new_G561_;
  assign new_G1023_ = ~new_G1689_ | ~new_G1692_;
  assign new_G1147_ = ~new_G1777_ | ~new_G1780_;
  assign new_G418_ = ~new_G416_ | ~new_G417_;
  assign new_G420_ = ~new_G1373_ | ~new_G1376_;
  assign new_G425_ = ~new_G423_ | ~new_G424_;
  assign new_G510_ = ~new_G508_ | ~new_G509_;
  assign new_G513_ = ~new_G511_ | ~new_G512_;
  assign new_G552_ = ~new_G546_;
  assign new_G1025_ = ~new_G1023_ | ~new_G1024_;
  assign new_G1149_ = ~new_G1147_ | ~new_G1148_;
  assign new_G419_ = ~new_G418_;
  assign new_G422_ = ~new_G420_ | ~new_G421_;
  assign new_G441_ = ~new_G425_ | ~new_G918_;
  assign new_G516_ = ~new_G510_;
  assign new_G725_ = ~new_G549_;
  assign new_G728_ = new_G549_;
  assign new_G1029_ = ~new_G1025_;
  assign new_G1153_ = ~new_G1149_;
  assign new_G433_ = ~new_G419_ | ~new_G918_;
  assign new_G437_ = ~new_G422_ | ~new_G918_;
  assign new_G663_ = ~new_G513_;
  assign new_G666_ = new_G513_;
  assign new_G731_ = new_G719_ & new_G725_;
  assign new_G746_ = new_G722_ & new_G725_;
  assign new_G756_ = new_G719_ & new_G728_;
  assign new_G770_ = new_G722_ & new_G728_;
  assign new_G1461_ = new_G441_;
  assign new_G1469_ = new_G441_;
  assign new_G1413_ = new_G433_;
  assign new_G1421_ = new_G433_;
  assign new_G1445_ = new_G437_;
  assign new_G1453_ = new_G437_;
  assign new_G532_ = ~new_G1469_ | ~new_G1472_;
  assign new_G1473_ = ~new_G1469_;
  assign new_G535_ = ~new_G1461_ | ~new_G1464_;
  assign new_G1465_ = ~new_G1461_;
  assign new_G495_ = ~new_G1421_ | ~new_G1424_;
  assign new_G1425_ = ~new_G1421_;
  assign new_G498_ = ~new_G1413_ | ~new_G1416_;
  assign new_G1417_ = ~new_G1413_;
  assign new_G520_ = ~new_G1453_ | ~new_G1456_;
  assign new_G1457_ = ~new_G1453_;
  assign new_G523_ = ~new_G1445_ | ~new_G1448_;
  assign new_G1449_ = ~new_G1445_;
  assign new_G533_ = ~new_G1466_ | ~new_G1473_;
  assign new_G536_ = ~new_G1458_ | ~new_G1465_;
  assign new_G496_ = ~new_G1418_ | ~new_G1425_;
  assign new_G499_ = ~new_G1410_ | ~new_G1417_;
  assign new_G521_ = ~new_G1450_ | ~new_G1457_;
  assign new_G524_ = ~new_G1442_ | ~new_G1449_;
  assign new_G534_ = ~new_G532_ | ~new_G533_;
  assign new_G537_ = ~new_G535_ | ~new_G536_;
  assign new_G497_ = ~new_G495_ | ~new_G496_;
  assign new_G500_ = ~new_G498_ | ~new_G499_;
  assign new_G522_ = ~new_G520_ | ~new_G521_;
  assign new_G525_ = ~new_G523_ | ~new_G524_;
  assign new_G540_ = ~new_G534_;
  assign new_G503_ = ~new_G497_;
  assign new_G528_ = ~new_G522_;
  assign new_G669_ = ~new_G537_;
  assign new_G672_ = new_G537_;
  assign new_G569_ = ~new_G500_;
  assign new_G588_ = new_G566_ & new_G500_;
  assign new_G618_ = ~new_G525_;
  assign new_G639_ = new_G615_ & new_G525_;
  assign new_G867_ = ~new_G487_ | ~new_G503_ | ~new_G528_ | ~new_G482_ | ~new_G540_ | ~new_G552_ | ~new_G516_ | ~new_G564_;
  assign new_G588a_ = new_G588_;
  assign new_G588b_ = new_G588_;
  assign new_G639a_ = new_G639_;
  assign new_G639b_ = new_G639_;
  assign new_G675_ = new_G663_ & new_G669_;
  assign new_G688_ = new_G666_ & new_G669_;
  assign new_G696_ = new_G663_ & new_G672_;
  assign new_G710_ = new_G666_ & new_G672_;
  assign new_G73_ = new_G932_ & new_G932_ & new_G949_ & new_G867_;
  assign new_G572_ = new_G565_ & new_G569_;
  assign new_G573_ = new_G566_ & new_G569_;
  assign new_G621_ = new_G614_ & new_G618_;
  assign new_G622_ = new_G615_ & new_G618_;
  assign new_G776_ = ~new_G958_ | ~new_G731_ | ~new_G696_ | ~new_G588a_ | ~new_G639a_;
  assign new_G780_ = ~new_G958_ | ~new_G756_ | ~new_G675_ | ~new_G588a_ | ~new_G639a_;
  assign new_G784_ = ~new_G958_ | ~new_G746_ | ~new_G675_ | ~new_G588a_ | ~new_G639a_;
  assign new_G788_ = ~new_G958_ | ~new_G731_ | ~new_G688_ | ~new_G588a_ | ~new_G639a_;
  assign new_G812_ = ~new_G969_ | ~new_G746_ | ~new_G710_ | ~new_G588b_ | ~new_G639a_;
  assign new_G832_ = ~new_G969_ | ~new_G770_ | ~new_G696_ | ~new_G588b_ | ~new_G639b_;
  assign new_G836_ = ~new_G969_ | ~new_G756_ | ~new_G710_ | ~new_G588b_ | ~new_G639b_;
  assign new_G1509_ = new_G958_ & new_G731_ & new_G696_ & new_G588a_ & new_G639a_;
  assign new_G1517_ = new_G958_ & new_G756_ & new_G675_ & new_G588a_ & new_G639a_;
  assign new_G1525_ = new_G958_ & new_G746_ & new_G675_ & new_G588a_ & new_G639a_;
  assign new_G1533_ = new_G958_ & new_G731_ & new_G688_ & new_G588a_ & new_G639a_;
  assign new_G1581_ = new_G969_ & new_G746_ & new_G710_ & new_G588b_ & new_G639a_;
  assign new_G1621_ = new_G969_ & new_G770_ & new_G696_ & new_G588b_ & new_G639b_;
  assign new_G1629_ = new_G969_ & new_G756_ & new_G710_ & new_G588b_ & new_G639b_;
  assign new_G792_ = ~new_G958_ | ~new_G756_ | ~new_G696_ | ~new_G588a_ | ~new_G622_;
  assign new_G796_ = ~new_G958_ | ~new_G746_ | ~new_G696_ | ~new_G588b_ | ~new_G622_;
  assign new_G800_ = ~new_G958_ | ~new_G731_ | ~new_G710_ | ~new_G588b_ | ~new_G622_;
  assign new_G804_ = ~new_G958_ | ~new_G770_ | ~new_G675_ | ~new_G588b_ | ~new_G622_;
  assign new_G808_ = ~new_G969_ | ~new_G756_ | ~new_G688_ | ~new_G588b_ | ~new_G622_;
  assign new_G816_ = ~new_G969_ | ~new_G756_ | ~new_G696_ | ~new_G573_ | ~new_G639b_;
  assign new_G820_ = ~new_G969_ | ~new_G746_ | ~new_G696_ | ~new_G573_ | ~new_G639b_;
  assign new_G824_ = ~new_G969_ | ~new_G731_ | ~new_G710_ | ~new_G573_ | ~new_G639b_;
  assign new_G828_ = ~new_G969_ | ~new_G756_ | ~new_G688_ | ~new_G573_ | ~new_G639b_;
  assign new_G871_ = ~new_G979_ | ~new_G731_ | ~new_G675_ | ~new_G588b_ | ~new_G622_;
  assign new_G873_ = ~new_G979_ | ~new_G731_ | ~new_G675_ | ~new_G573_ | ~new_G639b_;
  assign new_G875_ = ~new_G979_ | ~new_G731_ | ~new_G696_ | ~new_G573_ | ~new_G622_;
  assign new_G877_ = ~new_G979_ | ~new_G756_ | ~new_G675_ | ~new_G573_ | ~new_G622_;
  assign new_G879_ = ~new_G979_ | ~new_G746_ | ~new_G675_ | ~new_G573_ | ~new_G622_;
  assign new_G881_ = ~new_G979_ | ~new_G731_ | ~new_G688_ | ~new_G573_ | ~new_G622_;
  assign new_G883_ = ~new_G979_ | ~new_G731_ | ~new_G675_ | ~new_G573_ | ~new_G621_;
  assign new_G885_ = ~new_G979_ | ~new_G731_ | ~new_G675_ | ~new_G572_ | ~new_G622_;
  assign new_G1541_ = new_G958_ & new_G756_ & new_G696_ & new_G588a_ & new_G622_;
  assign new_G1549_ = new_G958_ & new_G746_ & new_G696_ & new_G588b_ & new_G622_;
  assign new_G1557_ = new_G958_ & new_G731_ & new_G710_ & new_G588b_ & new_G622_;
  assign new_G1565_ = new_G958_ & new_G770_ & new_G675_ & new_G588b_ & new_G622_;
  assign new_G1573_ = new_G969_ & new_G756_ & new_G688_ & new_G588b_ & new_G622_;
  assign new_G1589_ = new_G969_ & new_G756_ & new_G696_ & new_G573_ & new_G639b_;
  assign new_G1597_ = new_G969_ & new_G746_ & new_G696_ & new_G573_ & new_G639b_;
  assign new_G1605_ = new_G969_ & new_G731_ & new_G710_ & new_G573_ & new_G639b_;
  assign new_G1613_ = new_G969_ & new_G756_ & new_G688_ & new_G573_ & new_G639b_;
  assign new_G1_ = ~new_G1509_ | ~new_G1512_;
  assign new_G1513_ = ~new_G1509_;
  assign new_G4_ = ~new_G1517_ | ~new_G1520_;
  assign new_G1521_ = ~new_G1517_;
  assign new_G7_ = ~new_G1525_ | ~new_G1528_;
  assign new_G1529_ = ~new_G1525_;
  assign new_G10_ = ~new_G1533_ | ~new_G1536_;
  assign new_G1537_ = ~new_G1533_;
  assign new_G28_ = ~new_G1581_ | ~new_G1584_;
  assign new_G1585_ = ~new_G1581_;
  assign new_G43_ = ~new_G1621_ | ~new_G1624_;
  assign new_G1625_ = ~new_G1621_;
  assign new_G46_ = ~new_G1629_ | ~new_G1632_;
  assign new_G1633_ = ~new_G1629_;
  assign new_G886_ = new_G885_ & new_G883_ & new_G881_ & new_G879_ & new_G877_ & new_G875_ & new_G871_ & new_G873_;
  assign new_G2_ = ~new_G1506_ | ~new_G1513_;
  assign new_G5_ = ~new_G1514_ | ~new_G1521_;
  assign new_G8_ = ~new_G1522_ | ~new_G1529_;
  assign new_G11_ = ~new_G1530_ | ~new_G1537_;
  assign new_G13_ = ~new_G1541_ | ~new_G1544_;
  assign new_G1545_ = ~new_G1541_;
  assign new_G16_ = ~new_G1549_ | ~new_G1552_;
  assign new_G1553_ = ~new_G1549_;
  assign new_G19_ = ~new_G1557_ | ~new_G1560_;
  assign new_G1561_ = ~new_G1557_;
  assign new_G22_ = ~new_G1565_ | ~new_G1568_;
  assign new_G1569_ = ~new_G1565_;
  assign new_G25_ = ~new_G1573_ | ~new_G1576_;
  assign new_G1577_ = ~new_G1573_;
  assign new_G29_ = ~new_G1578_ | ~new_G1585_;
  assign new_G31_ = ~new_G1589_ | ~new_G1592_;
  assign new_G1593_ = ~new_G1589_;
  assign new_G34_ = ~new_G1597_ | ~new_G1600_;
  assign new_G1601_ = ~new_G1597_;
  assign new_G37_ = ~new_G1605_ | ~new_G1608_;
  assign new_G1609_ = ~new_G1605_;
  assign new_G40_ = ~new_G1613_ | ~new_G1616_;
  assign new_G1617_ = ~new_G1613_;
  assign new_G44_ = ~new_G1618_ | ~new_G1625_;
  assign new_G47_ = ~new_G1626_ | ~new_G1633_;
  assign new_G857_ = ~new_G804_ | ~new_G800_ | ~new_G796_ | ~new_G792_ | ~new_G788_ | ~new_G784_ | ~new_G776_ | ~new_G780_;
  assign new_G860_ = ~new_G836_ | ~new_G832_ | ~new_G828_ | ~new_G824_ | ~new_G820_ | ~new_G816_ | ~new_G808_ | ~new_G812_;
  assign new_G863_ = new_G804_ & new_G800_ & new_G796_ & new_G792_ & new_G788_ & new_G784_ & new_G776_ & new_G780_;
  assign new_G865_ = new_G836_ & new_G832_ & new_G828_ & new_G824_ & new_G820_ & new_G816_ & new_G808_ & new_G812_;
  assign G3 = ~new_G1_ | ~new_G2_;
  assign G6 = ~new_G4_ | ~new_G5_;
  assign G9 = ~new_G7_ | ~new_G8_;
  assign G12 = ~new_G10_ | ~new_G11_;
  assign new_G14_ = ~new_G1538_ | ~new_G1545_;
  assign new_G17_ = ~new_G1546_ | ~new_G1553_;
  assign new_G20_ = ~new_G1554_ | ~new_G1561_;
  assign new_G23_ = ~new_G1562_ | ~new_G1569_;
  assign new_G26_ = ~new_G1570_ | ~new_G1577_;
  assign G30 = ~new_G28_ | ~new_G29_;
  assign new_G32_ = ~new_G1586_ | ~new_G1593_;
  assign new_G35_ = ~new_G1594_ | ~new_G1601_;
  assign new_G38_ = ~new_G1602_ | ~new_G1609_;
  assign new_G41_ = ~new_G1610_ | ~new_G1617_;
  assign G45 = ~new_G43_ | ~new_G44_;
  assign G48 = ~new_G46_ | ~new_G47_;
  assign new_G1913_ = new_G857_ & new_G859_;
  assign new_G1921_ = new_G860_ & new_G862_;
  assign G15 = ~new_G13_ | ~new_G14_;
  assign G18 = ~new_G16_ | ~new_G17_;
  assign G21 = ~new_G19_ | ~new_G20_;
  assign G24 = ~new_G22_ | ~new_G23_;
  assign G27 = ~new_G25_ | ~new_G26_;
  assign G33 = ~new_G31_ | ~new_G32_;
  assign G36 = ~new_G34_ | ~new_G35_;
  assign G39 = ~new_G37_ | ~new_G38_;
  assign G42 = ~new_G40_ | ~new_G41_;
  assign new_G887_ = new_G886_ & new_G863_ & new_G865_;
  assign new_G462_ = ~new_G863_ | ~new_G865_;
  assign new_G74_ = new_G887_ & G952 & new_G949_ & new_G867_;
  assign new_G1637_ = ~new_G1913_ | ~new_G1916_;
  assign new_G1917_ = ~new_G1913_;
  assign new_G1647_ = ~new_G1921_ | ~new_G1924_;
  assign new_G1925_ = ~new_G1921_;
  assign G75 = ~new_G73_ & ~new_G74_;
  assign new_G1020_ = new_G462_ & new_G457_ & new_G911_;
  assign new_G1144_ = new_G462_ & G469 & new_G911_;
  assign new_G1386_ = new_G462_ & G475 & new_G911_;
  assign new_G1394_ = new_G462_ & G478 & new_G911_;
  assign new_G1402_ = new_G462_ & new_G459_ & new_G911_;
  assign new_G1638_ = ~new_G1910_ | ~new_G1917_;
  assign new_G1648_ = ~new_G1918_ | ~new_G1925_;
  assign new_G1806_ = new_G462_ & G472 & new_G911_;
  assign new_G1639_ = ~new_G1637_ | ~new_G1638_;
  assign new_G1649_ = ~new_G1647_ | ~new_G1648_;
  assign new_G287_ = ~new_G1020_ | ~new_G1029_;
  assign new_G350_ = ~new_G1144_ | ~new_G1153_;
  assign new_G427_ = ~new_G1386_ | ~new_G1393_;
  assign new_G429_ = ~new_G1394_ | ~new_G1401_;
  assign new_G431_ = ~new_G1402_ | ~new_G1409_;
  assign new_G1028_ = ~new_G1020_;
  assign new_G1152_ = ~new_G1144_;
  assign new_G1392_ = ~new_G1386_;
  assign new_G1400_ = ~new_G1394_;
  assign new_G1408_ = ~new_G1402_;
  assign new_G1812_ = ~new_G1806_;
  assign new_G1216_ = ~new_G1806_ | ~new_G1813_;
  assign new_G286_ = ~new_G1025_ | ~new_G1028_;
  assign new_G349_ = ~new_G1149_ | ~new_G1152_;
  assign new_G426_ = ~new_G1389_ | ~new_G1392_;
  assign new_G428_ = ~new_G1397_ | ~new_G1400_;
  assign new_G430_ = ~new_G1405_ | ~new_G1408_;
  assign new_G67_ = ~new_G1639_ | ~new_G1642_;
  assign new_G1643_ = ~new_G1639_;
  assign new_G70_ = ~new_G1649_ | ~new_G1652_;
  assign new_G1653_ = ~new_G1649_;
  assign new_G1215_ = ~new_G1809_ | ~new_G1812_;
  assign new_G49_ = ~new_G286_ | ~new_G287_;
  assign new_G53_ = ~new_G349_ | ~new_G350_;
  assign new_G59_ = ~new_G426_ | ~new_G427_;
  assign new_G61_ = ~new_G428_ | ~new_G429_;
  assign new_G65_ = ~new_G430_ | ~new_G431_;
  assign new_G68_ = ~new_G1634_ | ~new_G1643_;
  assign new_G71_ = ~new_G1644_ | ~new_G1653_;
  assign new_G1217_ = ~new_G1215_ | ~new_G1216_;
  assign G51 = new_G49_ & new_G50_;
  assign G54 = new_G52_ & new_G53_;
  assign G60 = new_G58_ & new_G59_;
  assign G63 = new_G61_ & new_G62_;
  assign G66 = new_G64_ & new_G65_;
  assign G69 = ~new_G67_ | ~new_G68_;
  assign G72 = ~new_G70_ | ~new_G71_;
  assign new_G375_ = ~new_G1217_ | ~new_G1220_;
  assign new_G1221_ = ~new_G1217_;
  assign new_G376_ = ~new_G1212_ | ~new_G1221_;
  assign new_G55_ = ~new_G375_ | ~new_G376_;
  assign G57 = new_G55_ & new_G56_;
endmodule


