// NOR_NOT mapped module c1908

module c1908 (
  input  G101    ,
  input  G104    ,
  input  G107    ,
  input  G110    ,
  input  G113    ,
  input  G116    ,
  input  G119    ,
  input  G122    ,
  input  G125    ,
  input  G128    ,
  input  G131    ,
  input  G134    ,
  input  G137    ,
  input  G140    ,
  input  G143    ,
  input  G146    ,
  input  G210    ,
  input  G214    ,
  input  G217    ,
  input  G221    ,
  input  G224    ,
  input  G227    ,
  input  G234    ,
  input  G237    ,
  input  G469    ,
  input  G472    ,
  input  G475    ,
  input  G478    ,
  input  G898    ,
  input  G900    ,
  input  G902    ,
  input  G952    ,
  input  G953    ,
  output G3      ,
  output G6      ,
  output G9      ,
  output G12     ,
  output G30     ,
  output G45     ,
  output G48     ,
  output G15     ,
  output G18     ,
  output G21     ,
  output G24     ,
  output G27     ,
  output G33     ,
  output G36     ,
  output G39     ,
  output G42     ,
  output G75     ,
  output G51     ,
  output G54     ,
  output G60     ,
  output G63     ,
  output G66     ,
  output G69     ,
  output G72     ,
  output G57     );

  wire wr_26;
  wire wr_27;
  wire wr_28;
  wire wr_29;
  wire wr_30;
  wire wr_31;
  wire wr_32;
  wire wr_33;
  wire wr_34;
  wire wr_35;
  wire wr_36;
  wire wr_37;
  wire wr_38;
  wire wr_39;
  wire wr_40;
  wire wr_41;
  wire wr_42;
  wire wr_43;
  wire wr_44;
  wire wr_45;
  wire wr_46;
  wire wr_47;
  wire wr_48;
  wire wr_49;
  wire wr_50;
  wire wr_51;
  wire wr_52;
  wire wr_53;
  wire wr_54;
  wire wr_55;
  wire wr_56;
  wire wr_57;
  wire wr_58;
  wire wr_59;
  wire wr_60;
  wire wr_61;
  wire wr_62;
  wire wr_63;
  wire wr_64;
  wire wr_65;
  wire wr_66;
  wire wr_67;
  wire wr_68;
  wire wr_69;
  wire wr_70;
  wire wr_71;
  wire wr_72;
  wire wr_73;
  wire wr_74;
  wire wr_75;
  wire wr_76;
  wire wr_77;
  wire wr_78;
  wire wr_79;
  wire wr_80;
  wire wr_81;
  wire wr_82;
  wire wr_83;
  wire wr_84;
  wire wr_85;
  wire wr_86;
  wire wr_87;
  wire wr_88;
  wire wr_89;
  wire wr_90;
  wire wr_91;
  wire wr_92;
  wire wr_93;
  wire wr_94;
  wire wr_95;
  wire wr_96;
  wire wr_97;
  wire wr_98;
  wire wr_99;
  wire wr_100;
  wire wr_101;
  wire wr_102;
  wire wr_103;
  wire wr_104;
  wire wr_105;
  wire wr_106;
  wire wr_107;
  wire wr_108;
  wire wr_109;
  wire wr_110;
  wire wr_111;
  wire wr_112;
  wire wr_113;
  wire wr_114;
  wire wr_115;
  wire wr_116;
  wire wr_117;
  wire wr_118;
  wire wr_119;
  wire wr_120;
  wire wr_121;
  wire wr_122;
  wire wr_123;
  wire wr_124;
  wire wr_125;
  wire wr_126;
  wire wr_127;
  wire wr_128;
  wire wr_129;
  wire wr_130;
  wire wr_131;
  wire wr_132;
  wire wr_133;
  wire wr_134;
  wire wr_135;
  wire wr_136;
  wire wr_137;
  wire wr_138;
  wire wr_139;
  wire wr_140;
  wire wr_141;
  wire wr_142;
  wire wr_143;
  wire wr_144;
  wire wr_145;
  wire wr_146;
  wire wr_147;
  wire wr_148;
  wire wr_149;
  wire wr_150;
  wire wr_151;
  wire wr_152;
  wire wr_153;
  wire wr_154;
  wire wr_155;
  wire wr_156;
  wire wr_157;
  wire wr_158;
  wire wr_159;
  wire wr_160;
  wire wr_161;
  wire wr_162;
  wire wr_163;
  wire wr_164;
  wire wr_165;
  wire wr_166;
  wire wr_167;
  wire wr_168;
  wire wr_169;
  wire wr_170;
  wire wr_171;
  wire wr_172;
  wire wr_173;
  wire wr_174;
  wire wr_175;
  wire wr_176;
  wire wr_177;
  wire wr_178;
  wire wr_179;
  wire wr_180;
  wire wr_181;
  wire wr_182;
  wire wr_183;
  wire wr_184;
  wire wr_185;
  wire wr_186;
  wire wr_187;
  wire wr_188;
  wire wr_189;
  wire wr_190;
  wire wr_191;
  wire wr_192;
  wire wr_193;
  wire wr_194;
  wire wr_195;
  wire wr_196;
  wire wr_197;
  wire wr_198;
  wire wr_199;
  wire wr_200;
  wire wr_201;
  wire wr_202;
  wire wr_203;
  wire wr_204;
  wire wr_205;
  wire wr_206;
  wire wr_207;
  wire wr_208;
  wire wr_209;
  wire wr_210;
  wire wr_211;
  wire wr_212;
  wire wr_213;
  wire wr_214;
  wire wr_215;
  wire wr_216;
  wire wr_217;
  wire wr_218;
  wire wr_219;
  wire wr_220;
  wire wr_221;
  wire wr_222;
  wire wr_223;
  wire wr_224;
  wire wr_225;
  wire wr_226;
  wire wr_227;
  wire wr_228;
  wire wr_229;
  wire wr_230;
  wire wr_231;
  wire wr_232;
  wire wr_233;
  wire wr_234;
  wire wr_235;
  wire wr_236;
  wire wr_237;
  wire wr_238;
  wire wr_239;
  wire wr_240;
  wire wr_241;
  wire wr_242;
  wire wr_243;
  wire wr_244;
  wire wr_245;
  wire wr_246;
  wire wr_247;
  wire wr_248;
  wire wr_249;
  wire wr_250;
  wire wr_251;
  wire wr_252;
  wire wr_253;
  wire wr_254;
  wire wr_255;
  wire wr_256;
  wire wr_257;
  wire wr_258;
  wire wr_259;
  wire wr_260;
  wire wr_261;
  wire wr_262;
  wire wr_263;
  wire wr_264;
  wire wr_265;
  wire wr_266;
  wire wr_267;
  wire wr_268;
  wire wr_269;
  wire wr_270;
  wire wr_271;
  wire wr_272;
  wire wr_273;
  wire wr_274;
  wire wr_275;
  wire wr_276;
  wire wr_277;
  wire wr_278;
  wire wr_279;
  wire wr_280;
  wire wr_281;
  wire wr_282;
  wire wr_283;
  wire wr_284;
  wire wr_285;
  wire wr_286;
  wire wr_287;
  wire wr_288;
  wire wr_289;
  wire wr_290;
  wire wr_291;
  wire wr_292;
  wire wr_293;
  wire wr_294;
  wire wr_295;
  wire wr_296;
  wire wr_297;
  wire wr_298;
  wire wr_299;
  wire wr_300;
  wire wr_301;
  wire wr_302;
  wire wr_303;
  wire wr_304;
  wire wr_305;
  wire wr_306;
  wire wr_307;
  wire wr_308;
  wire wr_309;
  wire wr_310;
  wire wr_311;
  wire wr_312;
  wire wr_313;
  wire wr_314;
  wire wr_315;
  wire wr_316;
  wire wr_317;
  wire wr_318;
  wire wr_319;
  wire wr_320;
  wire wr_321;
  wire wr_322;
  wire wr_323;
  wire wr_324;
  wire wr_325;
  wire wr_326;
  wire wr_327;
  wire wr_328;
  wire wr_329;
  wire wr_330;
  wire wr_331;
  wire wr_332;
  wire wr_333;
  wire wr_334;
  wire wr_335;
  wire wr_336;
  wire wr_337;
  wire wr_338;
  wire wr_339;
  wire wr_340;
  wire wr_341;
  wire wr_342;
  wire wr_343;
  wire wr_344;
  wire wr_345;
  wire wr_346;
  wire wr_347;
  wire wr_348;
  wire wr_349;
  wire wr_350;
  wire wr_351;
  wire wr_352;
  wire wr_353;
  wire wr_354;
  wire wr_355;
  wire wr_356;
  wire wr_357;
  wire wr_358;
  wire wr_359;
  wire wr_360;
  wire wr_361;
  wire wr_362;
  wire wr_363;
  wire wr_364;
  wire wr_365;
  wire wr_366;
  wire wr_367;
  wire wr_368;
  wire wr_369;
  wire wr_370;
  wire wr_371;
  wire wr_372;
  wire wr_373;
  wire wr_374;
  wire wr_375;
  wire wr_376;
  wire wr_377;
  wire wr_378;
  wire wr_379;
  wire wr_380;
  wire wr_381;
  wire wr_382;
  wire wr_383;
  wire wr_384;
  wire wr_385;
  wire wr_386;
  wire wr_387;
  wire wr_388;
  wire wr_389;
  wire wr_390;
  wire wr_391;
  wire wr_392;
  wire wr_393;
  wire wr_394;
  wire wr_395;
  wire wr_396;
  wire wr_397;
  wire wr_398;
  wire wr_399;
  wire wr_400;
  wire wr_401;
  wire wr_402;
  wire wr_403;
  wire wr_404;
  wire wr_405;
  wire wr_406;
  wire wr_407;
  wire wr_408;
  wire wr_409;
  wire wr_410;
  wire wr_411;
  wire wr_412;
  wire wr_413;
  wire wr_414;
  wire wr_415;
  wire wr_416;
  wire wr_417;
  wire wr_418;
  wire wr_419;
  wire wr_420;
  wire wr_421;
  wire wr_422;
  wire wr_423;
  wire wr_424;
  wire wr_425;
  wire wr_426;
  wire wr_427;
  wire wr_428;
  wire wr_429;
  wire wr_430;
  wire wr_431;
  wire wr_432;
  wire wr_433;
  wire wr_434;
  wire wr_435;
  wire wr_436;
  wire wr_437;
  wire wr_438;
  wire wr_439;
  wire wr_440;
  wire wr_441;
  wire wr_442;
  wire wr_443;
  wire wr_444;
  wire wr_445;
  wire wr_446;
  wire wr_447;
  wire wr_448;
  wire wr_449;
  wire wr_450;
  wire wr_451;
  wire wr_452;
  wire wr_453;
  wire wr_454;
  wire wr_455;
  wire wr_456;
  wire wr_457;
  wire wr_458;
  wire wr_459;
  wire wr_460;
  wire wr_461;
  wire wr_462;
  wire wr_463;
  wire wr_464;
  wire wr_465;
  wire wr_466;
  wire wr_467;
  wire wr_468;
  wire wr_469;
  wire wr_470;
  wire wr_471;
  wire wr_472;
  wire wr_473;
  wire wr_474;
  wire wr_475;
  wire wr_476;
  wire wr_477;
  wire wr_478;
  wire wr_479;
  wire wr_480;
  wire wr_481;
  wire wr_482;
  wire wr_483;
  wire wr_484;
  wire wr_485;
  wire wr_486;
  wire wr_487;
  wire wr_488;
  wire wr_489;
  wire wr_490;
  wire wr_491;
  wire wr_492;
  wire wr_493;
  wire wr_494;
  wire wr_495;
  wire wr_496;
  wire wr_497;
  wire wr_498;
  wire wr_499;
  wire wr_500;
  wire wr_501;
  wire wr_502;
  wire wr_503;
  wire wr_504;
  wire wr_505;
  wire wr_506;
  wire wr_507;
  wire wr_508;
  wire wr_509;
  wire wr_510;
  wire wr_511;
  wire wr_512;
  wire wr_513;
  wire wr_514;
  wire wr_515;
  wire wr_516;
  wire wr_517;
  wire wr_518;
  wire wr_519;
  wire wr_520;
  wire wr_521;
  wire wr_522;
  wire wr_523;
  wire wr_524;
  wire wr_525;
  wire wr_526;
  wire wr_527;
  wire wr_528;
  wire wr_529;
  wire wr_530;
  wire wr_531;
  wire wr_532;
  wire wr_533;
  wire wr_534;
  wire wr_535;
  wire wr_536;
  wire wr_537;
  wire wr_538;
  wire wr_539;
  wire wr_540;
  wire wr_541;
  wire wr_542;
  wire wr_543;
  wire wr_544;
  wire wr_545;
  wire wr_546;
  wire wr_547;
  wire wr_548;
  wire wr_549;
  wire wr_550;
  wire wr_551;
  wire wr_552;
  wire wr_553;
  wire wr_554;
  wire wr_555;
  wire wr_556;
  wire wr_557;
  wire wr_558;
  wire wr_559;
  wire wr_560;
  wire wr_561;
  wire wr_562;
  wire wr_563;
  wire wr_564;
  wire wr_565;
  wire wr_566;
  wire wr_567;
  wire wr_568;
  wire wr_569;
  wire wr_570;
  wire wr_571;
  wire wr_572;
  wire wr_573;
  wire wr_574;
  wire wr_575;
  wire wr_576;
  wire wr_577;
  wire wr_578;
  wire wr_579;
  wire wr_580;
  wire wr_581;
  wire wr_582;
  wire wr_583;
  wire wr_584;
  wire wr_585;
  wire wr_586;
  wire wr_587;
  wire wr_588;
  wire wr_589;
  wire wr_590;
  wire wr_591;
  wire wr_592;
  wire wr_593;
  wire wr_594;
  wire wr_595;
  wire wr_596;
  wire wr_597;
  wire wr_598;
  wire wr_599;
  wire wr_600;
  wire wr_601;
  wire wr_602;
  wire wr_603;
  wire wr_604;
  wire wr_605;
  wire wr_606;
  wire wr_607;
  wire wr_608;
  wire wr_609;
  wire wr_610;
  wire wr_611;
  wire wr_612;
  wire wr_613;
  wire wr_614;
  wire wr_615;
  wire wr_616;
  wire wr_617;
  wire wr_618;
  wire wr_619;
  wire wr_620;
  wire wr_621;
  wire wr_622;
  wire wr_623;
  wire wr_624;
  wire wr_625;
  wire wr_626;
  wire wr_627;
  wire wr_628;
  wire wr_629;
  wire wr_630;
  wire wr_631;
  wire wr_632;
  wire wr_633;
  wire wr_634;
  wire wr_635;
  wire wr_636;
  wire wr_637;
  wire wr_638;
  wire wr_639;
  wire wr_640;
  wire wr_641;
  wire wr_642;
  wire wr_643;
  wire wr_644;
  wire wr_645;
  wire wr_646;
  wire wr_647;
  wire wr_648;
  wire wr_649;
  wire wr_650;
  wire wr_651;
  wire wr_652;
  wire wr_653;
  wire wr_654;
  wire wr_655;
  wire wr_656;
  wire wr_657;
  wire wr_658;
  wire wr_659;
  wire wr_660;
  wire wr_661;
  wire wr_662;
  wire wr_663;
  wire wr_664;
  wire wr_665;
  wire wr_666;
  wire wr_667;
  wire wr_668;
  wire wr_669;
  wire wr_670;
  wire wr_671;
  wire wr_672;
  wire wr_673;
  wire wr_674;
  wire wr_675;
  wire wr_676;
  wire wr_677;
  wire wr_678;
  wire wr_679;
  wire wr_680;
  wire wr_681;
  wire wr_682;
  wire wr_683;

  not    g1( wr_26   ,           G221    );
  not    g2( wr_27   ,           G234    );
  not    g3( wr_31   ,           G140    );
  not    g4( wr_33   ,           G110    );
  not    g5( wr_36   ,           G227    );
  not    g6( wr_43   ,           G131    );
  not    g7( wr_44   ,           G134    );
  not    g8( wr_46   ,           G137    );
  not    g9( wr_53   ,           G128    );
  not   g10( wr_54   ,           G143    );
  not   g11( wr_56   ,           G146    );
  not   g12( wr_63   ,           G101    );
  not   g13( wr_64   ,           G104    );
  not   g14( wr_66   ,           G107    );
  not   g15( wr_95   ,           G214    );
  not   g16( wr_98   ,           G125    );
  not   g17( wr_102  ,           G224    );
  not   g18( wr_110  ,           G113    );
  not   g19( wr_111  ,           G116    );
  not   g20( wr_113  ,           G119    );
  not   g21( wr_125  ,           G122    );
  not   g22( wr_139  ,           G210    );
  not   g23( wr_180  ,           G217    );
  not   g24( wr_217  ,           G237    );
  not   g25( wr_216  ,           G953    );
  not   g26( wr_229  ,           G478    );
  not   g27( wr_263  ,           G475    );
  not   g28( wr_224  ,           G952    );
  not   g29( wr_188  ,           G472    );
  nor   g30( wr_96   , G902    , G237    );
  not   g31( wr_215  ,           G902    );
  not   g32( wr_30   ,           G469    );
  not   g33( wr_645  ,           G898    );
  not   g34( wr_665  ,           G900    );
  nor   g35( wr_493  , G953    , G952    );
  nor   g36( wr_32   , wr_31   , G110    );
  nor   g37( wr_34   , G140    , wr_33   );
  nor   g38( wr_37   , G953    , wr_36   );
  nor   g39( wr_45   , G137    , wr_44   );
  nor   g40( wr_47   , wr_46   , G134    );
  nor   g41( wr_55   , G146    , wr_54   );
  nor   g42( wr_57   , wr_56   , G143    );
  nor   g43( wr_65   , G107    , wr_64   );
  nor   g44( wr_67   , wr_66   , G104    );
  nor   g45( wr_103  , G953    , wr_102  );
  nor   g46( wr_112  , G119    , wr_111  );
  nor   g47( wr_114  , wr_113  , G116    );
  nor   g48( wr_124  , G122    , wr_33   );
  nor   g49( wr_126  , wr_125  , G110    );
  nor   g50( wr_148  , wr_31   , G125    );
  nor   g51( wr_149  , G140    , wr_98   );
  nor   g52( wr_156  , G128    , wr_113  );
  nor   g53( wr_157  , wr_53   , G119    );
  nor   g54( wr_167  , G953    , wr_26   );
  nor   g55( wr_189  , G953    , wr_139  );
  nor   g56( wr_230  , G122    , wr_111  );
  nor   g57( wr_231  , wr_125  , G116    );
  nor   g58( wr_237  , G143    , wr_53   );
  nor   g59( wr_238  , wr_54   , G128    );
  nor   g60( wr_249  , G953    , wr_180  );
  nor   g61( wr_264  , G953    , wr_95   );
  nor   g62( wr_279  , G122    , wr_110  );
  nor   g63( wr_280  , wr_125  , G113    );
  nor   g64( wr_218  , wr_217  , wr_27   );
  nor   g65( wr_28   , G902    , wr_27   );
  nor   g66( wr_140  , wr_96   , wr_139  );
  nor   g67( wr_97   , wr_96   , wr_95   );
  nor   g68( wr_639  , wr_216  , G898    );
  nor   g69( wr_655  , wr_216  , G900    );
  nor   g70( wr_646  , wr_645  , wr_102  );
  nor   g71( wr_666  , wr_665  , wr_36   );
  not   g72( wr_494  ,           wr_493  );
  nor   g73( wr_604  , wr_216  , G952    );
  nor   g74( wr_35   , wr_34   , wr_32   );
  nor   g75( wr_48   , wr_47   , wr_45   );
  nor   g76( wr_58   , wr_57   , wr_55   );
  nor   g77( wr_68   , wr_67   , wr_65   );
  not   g78( wr_106  ,           wr_103  );
  nor   g79( wr_115  , wr_114  , wr_112  );
  nor   g80( wr_127  , wr_126  , wr_124  );
  nor   g81( wr_150  , wr_149  , wr_148  );
  nor   g82( wr_158  , wr_157  , wr_156  );
  not   g83( wr_168  ,           wr_167  );
  not   g84( wr_190  ,           wr_189  );
  nor   g85( wr_232  , wr_231  , wr_230  );
  nor   g86( wr_239  , wr_238  , wr_237  );
  not   g87( wr_250  ,           wr_249  );
  not   g88( wr_265  ,           wr_264  );
  nor   g89( wr_281  , wr_280  , wr_279  );
  not   g90( wr_40   ,           wr_37   );
  nor   g91( wr_219  , wr_218  , wr_216  );
  nor   g92( wr_181  , wr_28   , wr_180  );
  nor   g93( wr_225  , wr_218  , wr_224  );
  not   g94( wr_141  ,           wr_140  );
  not   g95( wr_545  ,           wr_97   );
  nor   g96( wr_29   , wr_28   , wr_26   );
  nor   g97( wr_647  , wr_646  , wr_216  );
  nor   g98( wr_667  , wr_666  , wr_216  );
  nor   g99( wr_49   , wr_48   , wr_43   );
  not  g100( wr_50   ,           wr_48   );
  nor  g101( wr_59   , wr_58   , wr_53   );
  not  g102( wr_60   ,           wr_58   );
  nor  g103( wr_69   , wr_68   , wr_63   );
  not  g104( wr_70   ,           wr_68   );
  nor  g105( wr_116  , wr_115  , wr_110  );
  not  g106( wr_117  ,           wr_115  );
  not  g107( wr_130  ,           wr_127  );
  nor  g108( wr_151  , wr_150  , wr_56   );
  not  g109( wr_152  ,           wr_150  );
  nor  g110( wr_159  , wr_158  , wr_33   );
  not  g111( wr_160  ,           wr_158  );
  nor  g112( wr_169  , wr_168  , wr_27   );
  nor  g113( wr_191  , wr_190  , G237    );
  nor  g114( wr_233  , wr_232  , wr_66   );
  not  g115( wr_234  ,           wr_232  );
  nor  g116( wr_240  , wr_239  , wr_44   );
  not  g117( wr_241  ,           wr_239  );
  nor  g118( wr_251  , wr_250  , wr_27   );
  nor  g119( wr_266  , wr_265  , G237    );
  nor  g120( wr_282  , wr_281  , wr_64   );
  not  g121( wr_283  ,           wr_281  );
  not  g122( wr_39   ,           wr_35   );
  nor  g123( wr_38   , wr_37   , wr_35   );
  not  g124( wr_220  ,           wr_219  );
  not  g125( wr_182  ,           wr_181  );
  not  g126( wr_226  ,           wr_225  );
  not  g127( wr_551  ,           wr_29   );
  not  g128( wr_650  ,           wr_647  );
  not  g129( wr_670  ,           wr_667  );
  nor  g130( wr_51   , wr_50   , G131    );
  nor  g131( wr_61   , wr_60   , G128    );
  nor  g132( wr_71   , wr_70   , G101    );
  nor  g133( wr_118  , wr_117  , G113    );
  nor  g134( wr_153  , wr_152  , G146    );
  nor  g135( wr_161  , wr_160  , G110    );
  not  g136( wr_170  ,           wr_169  );
  nor  g137( wr_172  , wr_169  , G137    );
  nor  g138( wr_192  , wr_191  , G101    );
  not  g139( wr_193  ,           wr_191  );
  nor  g140( wr_235  , wr_234  , G107    );
  nor  g141( wr_242  , wr_241  , G134    );
  not  g142( wr_254  ,           wr_251  );
  nor  g143( wr_267  , wr_266  , G143    );
  not  g144( wr_268  ,           wr_266  );
  nor  g145( wr_284  , wr_283  , G104    );
  nor  g146( wr_41   , wr_40   , wr_39   );
  nor  g147( wr_221  , wr_220  , G898    );
  nor  g148( wr_352  , wr_220  , G900    );
  nor  g149( wr_227  , wr_226  , G953    );
  nor  g150( wr_52   , wr_51   , wr_49   );
  nor  g151( wr_62   , wr_61   , wr_59   );
  nor  g152( wr_72   , wr_71   , wr_69   );
  nor  g153( wr_119  , wr_118  , wr_116  );
  nor  g154( wr_154  , wr_153  , wr_151  );
  nor  g155( wr_162  , wr_161  , wr_159  );
  nor  g156( wr_171  , wr_170  , wr_46   );
  nor  g157( wr_194  , wr_193  , wr_63   );
  nor  g158( wr_236  , wr_235  , wr_233  );
  nor  g159( wr_243  , wr_242  , wr_240  );
  nor  g160( wr_269  , wr_268  , wr_54   );
  nor  g161( wr_285  , wr_284  , wr_282  );
  nor  g162( wr_42   , wr_41   , wr_38   );
  not  g163( wr_222  ,           wr_221  );
  not  g164( wr_353  ,           wr_352  );
  not  g165( wr_510  ,           wr_227  );
  nor  g166( wr_73   , wr_72   , wr_62   );
  not  g167( wr_74   ,           wr_62   );
  not  g168( wr_75   ,           wr_72   );
  not  g169( wr_79   ,           wr_52   );
  nor  g170( wr_99   , wr_62   , wr_98   );
  not  g171( wr_120  ,           wr_119  );
  nor  g172( wr_122  , wr_119  , wr_72   );
  not  g173( wr_155  ,           wr_154  );
  not  g174( wr_164  ,           wr_162  );
  nor  g175( wr_173  , wr_172  , wr_171  );
  nor  g176( wr_195  , wr_194  , wr_192  );
  nor  g177( wr_198  , wr_62   , wr_52   );
  not  g178( wr_244  ,           wr_243  );
  not  g179( wr_246  ,           wr_236  );
  nor  g180( wr_270  , wr_269  , wr_267  );
  not  g181( wr_286  ,           wr_285  );
  not  g182( wr_84   ,           wr_42   );
  nor  g183( wr_223  , wr_222  , wr_215  );
  nor  g184( wr_354  , wr_353  , wr_215  );
  nor  g185( wr_76   , wr_75   , wr_74   );
  nor  g186( wr_100  , wr_74   , G125    );
  nor  g187( wr_121  , wr_120  , wr_75   );
  nor  g188( wr_163  , wr_162  , wr_155  );
  nor  g189( wr_165  , wr_164  , wr_154  );
  not  g190( wr_176  ,           wr_173  );
  not  g191( wr_196  ,           wr_195  );
  nor  g192( wr_197  , wr_74   , wr_79   );
  nor  g193( wr_245  , wr_244  , wr_236  );
  nor  g194( wr_247  , wr_243  , wr_246  );
  nor  g195( wr_271  , wr_270  , wr_43   );
  not  g196( wr_272  ,           wr_270  );
  nor  g197( wr_228  , wr_227  , wr_223  );
  nor  g198( wr_355  , wr_354  , wr_227  );
  nor  g199( wr_77   , wr_76   , wr_73   );
  nor  g200( wr_101  , wr_100  , wr_99   );
  nor  g201( wr_123  , wr_122  , wr_121  );
  nor  g202( wr_166  , wr_165  , wr_163  );
  nor  g203( wr_199  , wr_198  , wr_197  );
  nor  g204( wr_248  , wr_247  , wr_245  );
  nor  g205( wr_273  , wr_272  , G131    );
  nor  g206( wr_104  , wr_103  , wr_101  );
  not  g207( wr_105  ,           wr_101  );
  nor  g208( wr_128  , wr_127  , wr_123  );
  not  g209( wr_129  ,           wr_123  );
  not  g210( wr_175  ,           wr_166  );
  nor  g211( wr_200  , wr_199  , wr_119  );
  not  g212( wr_201  ,           wr_199  );
  nor  g213( wr_252  , wr_251  , wr_248  );
  not  g214( wr_253  ,           wr_248  );
  nor  g215( wr_274  , wr_273  , wr_271  );
  not  g216( wr_80   ,           wr_77   );
  nor  g217( wr_174  , wr_173  , wr_166  );
  nor  g218( wr_78   , wr_77   , wr_52   );
  nor  g219( wr_656  , wr_199  , wr_150  );
  nor  g220( wr_107  , wr_106  , wr_105  );
  nor  g221( wr_131  , wr_130  , wr_129  );
  nor  g222( wr_202  , wr_201  , wr_120  );
  nor  g223( wr_255  , wr_254  , wr_253  );
  not  g224( wr_275  ,           wr_274  );
  nor  g225( wr_277  , wr_274  , wr_155  );
  nor  g226( wr_177  , wr_176  , wr_175  );
  nor  g227( wr_81   , wr_80   , wr_79   );
  nor  g228( wr_657  , wr_201  , wr_152  );
  nor  g229( wr_203  , wr_202  , wr_200  );
  nor  g230( wr_256  , wr_255  , wr_252  );
  nor  g231( wr_276  , wr_275  , wr_154  );
  nor  g232( wr_108  , wr_107  , wr_104  );
  nor  g233( wr_132  , wr_131  , wr_128  );
  nor  g234( wr_178  , wr_177  , wr_174  );
  nor  g235( wr_82   , wr_81   , wr_78   );
  nor  g236( wr_658  , wr_657  , wr_656  );
  not  g237( wr_205  ,           wr_203  );
  nor  g238( wr_278  , wr_277  , wr_276  );
  nor  g239( wr_204  , wr_203  , wr_196  );
  nor  g240( wr_257  , wr_256  , G902    );
  not  g241( wr_109  ,           wr_108  );
  not  g242( wr_133  ,           wr_132  );
  nor  g243( wr_135  , wr_132  , wr_108  );
  nor  g244( wr_179  , wr_178  , G902    );
  not  g245( wr_85   ,           wr_82   );
  nor  g246( wr_83   , wr_82   , wr_42   );
  not  g247( wr_659  ,           wr_658  );
  not  g248( wr_625  ,           wr_256  );
  not  g249( wr_633  ,           wr_178  );
  nor  g250( wr_287  , wr_286  , wr_278  );
  not  g251( wr_288  ,           wr_278  );
  nor  g252( wr_206  , wr_205  , wr_195  );
  not  g253( wr_259  ,           wr_257  );
  nor  g254( wr_134  , wr_133  , wr_109  );
  nor  g255( wr_258  , wr_257  , wr_229  );
  not  g256( wr_184  ,           wr_179  );
  nor  g257( wr_86   , wr_85   , wr_84   );
  nor  g258( wr_183  , wr_182  , wr_179  );
  nor  g259( wr_640  , wr_639  , wr_133  );
  nor  g260( wr_660  , wr_659  , wr_655  );
  nor  g261( wr_592  , wr_133  , wr_108  );
  nor  g262( wr_593  , wr_132  , wr_109  );
  nor  g263( wr_289  , wr_285  , wr_288  );
  nor  g264( wr_207  , wr_206  , wr_204  );
  nor  g265( wr_260  , wr_259  , G478    );
  nor  g266( wr_136  , wr_135  , wr_134  );
  nor  g267( wr_185  , wr_181  , wr_184  );
  nor  g268( wr_87   , wr_86   , wr_83   );
  not  g269( wr_642  ,           wr_640  );
  not  g270( wr_662  ,           wr_660  );
  nor  g271( wr_594  , wr_593  , wr_592  );
  nor  g272( wr_290  , wr_289  , wr_287  );
  nor  g273( wr_208  , wr_207  , G902    );
  nor  g274( wr_261  , wr_260  , wr_258  );
  not  g275( wr_137  ,           wr_136  );
  nor  g276( wr_186  , wr_185  , wr_183  );
  nor  g277( wr_88   , wr_87   , G902    );
  not  g278( wr_600  ,           wr_594  );
  not  g279( wr_609  ,           wr_87   );
  nor  g280( wr_291  , wr_290  , G902    );
  not  g281( wr_210  ,           wr_208  );
  nor  g282( wr_209  , wr_208  , wr_188  );
  not  g283( wr_262  ,           wr_261  );
  nor  g284( wr_138  , wr_137  , G902    );
  not  g285( wr_187  ,           wr_186  );
  not  g286( wr_90   ,           wr_88   );
  nor  g287( wr_89   , wr_88   , wr_30   );
  not  g288( wr_617  ,           wr_290  );
  not  g289( wr_293  ,           wr_291  );
  nor  g290( wr_292  , wr_291  , wr_263  );
  nor  g291( wr_211  , wr_210  , G472    );
  not  g292( wr_143  ,           wr_138  );
  nor  g293( wr_142  , wr_141  , wr_138  );
  nor  g294( wr_91   , wr_90   , G469    );
  nor  g295( wr_294  , wr_293  , G475    );
  nor  g296( wr_212  , wr_211  , wr_209  );
  nor  g297( wr_144  , wr_140  , wr_143  );
  nor  g298( wr_92   , wr_91   , wr_89   );
  nor  g299( wr_295  , wr_294  , wr_292  );
  not  g300( wr_310  ,           wr_212  );
  nor  g301( wr_213  , wr_212  , wr_187  );
  nor  g302( wr_350  , wr_212  , wr_186  );
  nor  g303( wr_145  , wr_144  , wr_142  );
  not  g304( wr_391  ,           wr_92   );
  nor  g305( wr_93   , wr_92   , wr_29   );
  not  g306( wr_296  ,           wr_295  );
  nor  g307( wr_313  , wr_295  , wr_262  );
  nor  g308( wr_367  , wr_295  , wr_261  );
  nor  g309( wr_311  , wr_310  , wr_187  );
  not  g310( wr_214  ,           wr_213  );
  not  g311( wr_351  ,           wr_350  );
  nor  g312( wr_146  , wr_145  , wr_97   );
  nor  g313( wr_339  , wr_310  , wr_186  );
  not  g314( wr_441  ,           wr_145  );
  nor  g315( wr_392  , wr_391  , wr_29   );
  not  g316( wr_94   ,           wr_93   );
  nor  g317( wr_552  , wr_391  , wr_551  );
  nor  g318( wr_297  , wr_296  , wr_262  );
  not  g319( wr_314  ,           wr_313  );
  not  g320( wr_368  ,           wr_367  );
  nor  g321( wr_326  , wr_296  , wr_261  );
  not  g322( wr_312  ,           wr_311  );
  not  g323( wr_147  ,           wr_146  );
  not  g324( wr_340  ,           wr_339  );
  nor  g325( wr_442  , wr_441  , wr_97   );
  nor  g326( wr_546  , wr_441  , wr_545  );
  not  g327( wr_393  ,           wr_392  );
  not  g328( wr_553  ,           wr_552  );
  nor  g329( wr_480  , wr_441  , wr_29   );
  not  g330( wr_298  ,           wr_297  );
  nor  g331( wr_369  , wr_368  , wr_355  );
  nor  g332( wr_380  , wr_355  , wr_314  );
  nor  g333( wr_421  , wr_368  , wr_228  );
  not  g334( wr_327  ,           wr_326  );
  nor  g335( wr_315  , wr_314  , wr_228  );
  not  g336( wr_443  ,           wr_442  );
  not  g337( wr_547  ,           wr_546  );
  nor  g338( wr_526  , wr_314  , wr_510  );
  not  g339( wr_481  ,           wr_480  );
  nor  g340( wr_299  , wr_298  , wr_228  );
  not  g341( wr_370  ,           wr_369  );
  not  g342( wr_381  ,           wr_380  );
  not  g343( wr_422  ,           wr_421  );
  nor  g344( wr_511  , wr_298  , wr_510  );
  nor  g345( wr_328  , wr_327  , wr_228  );
  nor  g346( wr_462  , wr_355  , wr_298  );
  not  g347( wr_316  ,           wr_315  );
  nor  g348( wr_533  , wr_327  , wr_510  );
  nor  g349( wr_356  , wr_355  , wr_327  );
  not  g350( wr_527  ,           wr_526  );
  nor  g351( wr_482  , wr_481  , wr_391  );
  not  g352( wr_300  ,           wr_299  );
  nor  g353( wr_371  , wr_370  , wr_214  );
  nor  g354( wr_382  , wr_381  , wr_351  );
  nor  g355( wr_423  , wr_422  , wr_312  );
  not  g356( wr_512  ,           wr_511  );
  not  g357( wr_329  ,           wr_328  );
  nor  g358( wr_432  , wr_381  , wr_340  );
  not  g359( wr_463  ,           wr_462  );
  nor  g360( wr_394  , wr_316  , wr_214  );
  not  g361( wr_534  ,           wr_533  );
  not  g362( wr_357  ,           wr_356  );
  nor  g363( wr_528  , wr_527  , wr_312  );
  nor  g364( wr_444  , wr_381  , wr_214  );
  nor  g365( wr_317  , wr_316  , wr_312  );
  not  g366( wr_483  ,           wr_482  );
  nor  g367( wr_412  , wr_351  , wr_300  );
  not  g368( wr_372  ,           wr_371  );
  not  g369( wr_383  ,           wr_382  );
  not  g370( wr_424  ,           wr_423  );
  nor  g371( wr_513  , wr_512  , wr_312  );
  nor  g372( wr_403  , wr_329  , wr_214  );
  not  g373( wr_433  ,           wr_432  );
  nor  g374( wr_540  , wr_512  , wr_340  );
  nor  g375( wr_464  , wr_463  , wr_351  );
  not  g376( wr_395  ,           wr_394  );
  nor  g377( wr_535  , wr_534  , wr_312  );
  nor  g378( wr_341  , wr_340  , wr_300  );
  nor  g379( wr_453  , wr_357  , wr_214  );
  nor  g380( wr_330  , wr_329  , wr_312  );
  not  g381( wr_529  ,           wr_528  );
  not  g382( wr_445  ,           wr_444  );
  nor  g383( wr_521  , wr_512  , wr_214  );
  nor  g384( wr_301  , wr_300  , wr_214  );
  nor  g385( wr_358  , wr_357  , wr_351  );
  not  g386( wr_318  ,           wr_317  );
  nor  g387( wr_484  , wr_483  , wr_97   );
  not  g388( wr_413  ,           wr_412  );
  nor  g389( wr_373  , wr_372  , wr_147  );
  nor  g390( wr_384  , wr_383  , wr_147  );
  nor  g391( wr_425  , wr_424  , wr_147  );
  not  g392( wr_514  ,           wr_513  );
  not  g393( wr_404  ,           wr_403  );
  nor  g394( wr_473  , wr_443  , wr_433  );
  not  g395( wr_541  ,           wr_540  );
  not  g396( wr_465  ,           wr_464  );
  nor  g397( wr_396  , wr_395  , wr_147  );
  not  g398( wr_536  ,           wr_535  );
  not  g399( wr_342  ,           wr_341  );
  not  g400( wr_454  ,           wr_453  );
  not  g401( wr_331  ,           wr_330  );
  nor  g402( wr_530  , wr_529  , wr_443  );
  nor  g403( wr_446  , wr_445  , wr_443  );
  not  g404( wr_522  ,           wr_521  );
  not  g405( wr_302  ,           wr_301  );
  nor  g406( wr_434  , wr_433  , wr_147  );
  not  g407( wr_359  ,           wr_358  );
  nor  g408( wr_319  , wr_318  , wr_147  );
  not  g409( wr_485  ,           wr_484  );
  nor  g410( wr_414  , wr_413  , wr_147  );
  not  g411( wr_374  ,           wr_373  );
  not  g412( wr_385  ,           wr_384  );
  not  g413( wr_426  ,           wr_425  );
  nor  g414( wr_515  , wr_514  , wr_443  );
  nor  g415( wr_548  , wr_547  , wr_514  );
  nor  g416( wr_405  , wr_404  , wr_147  );
  not  g417( wr_474  ,           wr_473  );
  nor  g418( wr_542  , wr_541  , wr_443  );
  nor  g419( wr_466  , wr_465  , wr_443  );
  not  g420( wr_397  ,           wr_396  );
  nor  g421( wr_537  , wr_536  , wr_443  );
  nor  g422( wr_343  , wr_342  , wr_147  );
  nor  g423( wr_455  , wr_454  , wr_443  );
  nor  g424( wr_332  , wr_331  , wr_147  );
  not  g425( wr_531  ,           wr_530  );
  not  g426( wr_447  ,           wr_446  );
  nor  g427( wr_523  , wr_522  , wr_443  );
  nor  g428( wr_303  , wr_302  , wr_147  );
  not  g429( wr_435  ,           wr_434  );
  nor  g430( wr_518  , wr_514  , wr_147  );
  nor  g431( wr_360  , wr_359  , wr_147  );
  not  g432( wr_320  ,           wr_319  );
  nor  g433( wr_486  , wr_485  , wr_310  );
  not  g434( wr_415  ,           wr_414  );
  nor  g435( wr_375  , wr_374  , wr_94   );
  nor  g436( wr_386  , wr_385  , wr_94   );
  nor  g437( wr_427  , wr_426  , wr_393  );
  not  g438( wr_516  ,           wr_515  );
  not  g439( wr_549  ,           wr_548  );
  not  g440( wr_406  ,           wr_405  );
  nor  g441( wr_475  , wr_474  , wr_94   );
  not  g442( wr_543  ,           wr_542  );
  not  g443( wr_467  ,           wr_466  );
  nor  g444( wr_398  , wr_397  , wr_393  );
  not  g445( wr_538  ,           wr_537  );
  not  g446( wr_344  ,           wr_343  );
  not  g447( wr_456  ,           wr_455  );
  not  g448( wr_333  ,           wr_332  );
  nor  g449( wr_532  , wr_531  , wr_393  );
  nor  g450( wr_448  , wr_447  , wr_94   );
  not  g451( wr_524  ,           wr_523  );
  not  g452( wr_304  ,           wr_303  );
  nor  g453( wr_436  , wr_435  , wr_393  );
  not  g454( wr_519  ,           wr_518  );
  not  g455( wr_361  ,           wr_360  );
  nor  g456( wr_321  , wr_320  , wr_94   );
  not  g457( wr_487  ,           wr_486  );
  nor  g458( wr_416  , wr_415  , wr_393  );
  nor  g459( wr_496  , wr_386  , wr_375  );
  nor  g460( wr_550  , wr_549  , wr_393  );
  nor  g461( wr_554  , wr_553  , wr_516  );
  nor  g462( wr_407  , wr_406  , wr_393  );
  nor  g463( wr_544  , wr_543  , wr_393  );
  nor  g464( wr_468  , wr_467  , wr_94   );
  nor  g465( wr_539  , wr_538  , wr_393  );
  nor  g466( wr_345  , wr_344  , wr_94   );
  nor  g467( wr_457  , wr_456  , wr_94   );
  nor  g468( wr_334  , wr_333  , wr_94   );
  nor  g469( wr_525  , wr_524  , wr_393  );
  nor  g470( wr_305  , wr_304  , wr_94   );
  nor  g471( wr_520  , wr_519  , wr_393  );
  nor  g472( wr_362  , wr_361  , wr_94   );
  nor  g473( wr_517  , wr_516  , wr_94   );
  nor  g474( wr_488  , wr_487  , wr_296  );
  not  g475( wr_322  ,           wr_321  );
  not  g476( wr_376  ,           wr_375  );
  not  g477( wr_387  ,           wr_386  );
  not  g478( wr_399  ,           wr_398  );
  not  g479( wr_428  ,           wr_427  );
  not  g480( wr_437  ,           wr_436  );
  not  g481( wr_449  ,           wr_448  );
  not  g482( wr_476  ,           wr_475  );
  nor  g483( wr_324  , wr_321  , wr_64   );
  nor  g484( wr_378  , wr_375  , wr_54   );
  nor  g485( wr_389  , wr_386  , wr_56   );
  nor  g486( wr_401  , wr_398  , wr_110  );
  nor  g487( wr_430  , wr_427  , wr_125  );
  nor  g488( wr_439  , wr_436  , wr_98   );
  nor  g489( wr_451  , wr_448  , wr_43   );
  nor  g490( wr_478  , wr_475  , wr_31   );
  nor  g491( wr_569  , wr_427  , wr_416  );
  not  g492( wr_497  ,           wr_496  );
  nor  g493( wr_555  , wr_554  , wr_550  );
  not  g494( wr_489  ,           wr_488  );
  not  g495( wr_306  ,           wr_305  );
  not  g496( wr_335  ,           wr_334  );
  not  g497( wr_346  ,           wr_345  );
  not  g498( wr_363  ,           wr_362  );
  not  g499( wr_408  ,           wr_407  );
  not  g500( wr_417  ,           wr_416  );
  not  g501( wr_458  ,           wr_457  );
  not  g502( wr_469  ,           wr_468  );
  nor  g503( wr_308  , wr_305  , wr_63   );
  nor  g504( wr_323  , wr_322  , G104    );
  nor  g505( wr_337  , wr_334  , wr_66   );
  nor  g506( wr_348  , wr_345  , wr_33   );
  nor  g507( wr_365  , wr_362  , wr_53   );
  nor  g508( wr_377  , wr_376  , G143    );
  nor  g509( wr_388  , wr_387  , G146    );
  nor  g510( wr_400  , wr_399  , G113    );
  nor  g511( wr_410  , wr_407  , wr_111  );
  nor  g512( wr_419  , wr_416  , wr_113  );
  nor  g513( wr_429  , wr_428  , G122    );
  nor  g514( wr_438  , wr_437  , G125    );
  nor  g515( wr_450  , wr_449  , G131    );
  nor  g516( wr_460  , wr_457  , wr_44   );
  nor  g517( wr_471  , wr_468  , wr_46   );
  nor  g518( wr_477  , wr_476  , G140    );
  not  g519( wr_570  ,           wr_569  );
  nor  g520( wr_498  , wr_497  , wr_475  );
  not  g521( wr_556  ,           wr_555  );
  nor  g522( wr_490  , wr_489  , wr_187  );
  nor  g523( wr_307  , wr_306  , G101    );
  nor  g524( wr_336  , wr_335  , G107    );
  nor  g525( wr_347  , wr_346  , G110    );
  nor  g526( wr_364  , wr_363  , G128    );
  nor  g527( wr_409  , wr_408  , G116    );
  nor  g528( wr_418  , wr_417  , G119    );
  nor  g529( wr_459  , wr_458  , G134    );
  nor  g530( wr_470  , wr_469  , G137    );
  nor  g531( wr_325  , wr_324  , wr_323  );
  nor  g532( wr_379  , wr_378  , wr_377  );
  nor  g533( wr_390  , wr_389  , wr_388  );
  nor  g534( wr_402  , wr_401  , wr_400  );
  nor  g535( wr_431  , wr_430  , wr_429  );
  nor  g536( wr_440  , wr_439  , wr_438  );
  nor  g537( wr_452  , wr_451  , wr_450  );
  nor  g538( wr_479  , wr_478  , wr_477  );
  nor  g539( wr_571  , wr_570  , wr_407  );
  not  g540( wr_499  ,           wr_498  );
  nor  g541( wr_557  , wr_556  , wr_544  );
  not  g542( wr_491  ,           wr_490  );
  nor  g543( wr_309  , wr_308  , wr_307  );
  nor  g544( wr_338  , wr_337  , wr_336  );
  nor  g545( wr_349  , wr_348  , wr_347  );
  nor  g546( wr_366  , wr_365  , wr_364  );
  nor  g547( wr_411  , wr_410  , wr_409  );
  nor  g548( wr_420  , wr_419  , wr_418  );
  nor  g549( wr_461  , wr_460  , wr_459  );
  nor  g550( wr_472  , wr_471  , wr_470  );
  not  g551( G6      ,           wr_325  );
  not  g552( G45     ,           wr_379  );
  not  g553( G48     ,           wr_390  );
  not  g554( G15     ,           wr_402  );
  not  g555( G24     ,           wr_431  );
  not  g556( G27     ,           wr_440  );
  not  g557( G33     ,           wr_452  );
  not  g558( G42     ,           wr_479  );
  not  g559( wr_572  ,           wr_571  );
  nor  g560( wr_500  , wr_499  , wr_468  );
  not  g561( wr_558  ,           wr_557  );
  nor  g562( wr_492  , wr_491  , wr_262  );
  not  g563( G3      ,           wr_309  );
  not  g564( G9      ,           wr_338  );
  not  g565( G12     ,           wr_349  );
  not  g566( G30     ,           wr_366  );
  not  g567( G18     ,           wr_411  );
  not  g568( G21     ,           wr_420  );
  not  g569( G36     ,           wr_461  );
  not  g570( G39     ,           wr_472  );
  nor  g571( wr_573  , wr_572  , wr_398  );
  not  g572( wr_501  ,           wr_500  );
  nor  g573( wr_559  , wr_558  , wr_539  );
  nor  g574( wr_495  , wr_494  , wr_492  );
  not  g575( wr_574  ,           wr_573  );
  nor  g576( wr_502  , wr_501  , wr_457  );
  not  g577( wr_560  ,           wr_559  );
  nor  g578( wr_575  , wr_574  , wr_345  );
  not  g579( wr_503  ,           wr_502  );
  nor  g580( wr_561  , wr_560  , wr_532  );
  not  g581( wr_576  ,           wr_575  );
  nor  g582( wr_504  , wr_503  , wr_448  );
  not  g583( wr_562  ,           wr_561  );
  nor  g584( wr_577  , wr_576  , wr_334  );
  not  g585( wr_505  ,           wr_504  );
  nor  g586( wr_563  , wr_562  , wr_525  );
  not  g587( wr_578  ,           wr_577  );
  nor  g588( wr_506  , wr_505  , wr_436  );
  not  g589( wr_564  ,           wr_563  );
  nor  g590( wr_579  , wr_578  , wr_305  );
  not  g591( wr_507  ,           wr_506  );
  nor  g592( wr_565  , wr_564  , wr_520  );
  not  g593( wr_580  ,           wr_579  );
  nor  g594( wr_508  , wr_507  , wr_362  );
  not  g595( wr_566  ,           wr_565  );
  nor  g596( wr_581  , wr_580  , wr_321  );
  not  g597( wr_509  ,           wr_508  );
  nor  g598( wr_567  , wr_566  , wr_517  );
  nor  g599( wr_653  , wr_508  , G953    );
  not  g600( wr_582  ,           wr_581  );
  not  g601( wr_568  ,           wr_567  );
  nor  g602( wr_637  , wr_581  , G953    );
  not  g603( wr_654  ,           wr_653  );
  nor  g604( wr_663  , wr_662  , wr_653  );
  nor  g605( wr_595  , wr_582  , wr_509  );
  nor  g606( wr_583  , wr_582  , wr_568  );
  not  g607( wr_638  ,           wr_637  );
  nor  g608( wr_643  , wr_642  , wr_637  );
  nor  g609( wr_661  , wr_660  , wr_654  );
  nor  g610( wr_673  , wr_595  , wr_188  );
  not  g611( wr_584  ,           wr_583  );
  nor  g612( wr_596  , wr_595  , wr_141  );
  nor  g613( wr_605  , wr_595  , wr_30   );
  nor  g614( wr_613  , wr_595  , wr_263  );
  nor  g615( wr_621  , wr_595  , wr_229  );
  nor  g616( wr_629  , wr_595  , wr_182  );
  nor  g617( wr_641  , wr_640  , wr_638  );
  nor  g618( wr_664  , wr_663  , wr_661  );
  not  g619( wr_674  ,           wr_673  );
  nor  g620( wr_585  , wr_584  , wr_509  );
  not  g621( wr_597  ,           wr_596  );
  not  g622( wr_606  ,           wr_605  );
  not  g623( wr_614  ,           wr_613  );
  not  g624( wr_622  ,           wr_621  );
  not  g625( wr_630  ,           wr_629  );
  nor  g626( wr_644  , wr_643  , wr_641  );
  not  g627( wr_669  ,           wr_664  );
  nor  g628( wr_668  , wr_667  , wr_664  );
  nor  g629( wr_675  , wr_674  , wr_215  );
  not  g630( wr_586  ,           wr_585  );
  nor  g631( wr_598  , wr_597  , wr_215  );
  nor  g632( wr_607  , wr_606  , wr_215  );
  nor  g633( wr_615  , wr_614  , wr_215  );
  nor  g634( wr_623  , wr_622  , wr_215  );
  nor  g635( wr_631  , wr_630  , wr_215  );
  not  g636( wr_649  ,           wr_644  );
  nor  g637( wr_648  , wr_647  , wr_644  );
  nor  g638( wr_671  , wr_670  , wr_669  );
  not  g639( wr_677  ,           wr_675  );
  nor  g640( wr_587  , wr_586  , wr_224  );
  nor  g641( wr_676  , wr_675  , wr_203  );
  not  g642( wr_601  ,           wr_598  );
  not  g643( wr_610  ,           wr_607  );
  not  g644( wr_618  ,           wr_615  );
  not  g645( wr_626  ,           wr_623  );
  not  g646( wr_634  ,           wr_631  );
  nor  g647( wr_599  , wr_598  , wr_594  );
  nor  g648( wr_608  , wr_607  , wr_87   );
  nor  g649( wr_616  , wr_615  , wr_290  );
  nor  g650( wr_624  , wr_623  , wr_256  );
  nor  g651( wr_632  , wr_631  , wr_178  );
  nor  g652( wr_651  , wr_650  , wr_649  );
  nor  g653( wr_672  , wr_671  , wr_668  );
  nor  g654( wr_678  , wr_677  , wr_205  );
  not  g655( wr_588  ,           wr_587  );
  nor  g656( wr_602  , wr_601  , wr_600  );
  nor  g657( wr_611  , wr_610  , wr_609  );
  nor  g658( wr_619  , wr_618  , wr_617  );
  nor  g659( wr_627  , wr_626  , wr_625  );
  nor  g660( wr_635  , wr_634  , wr_633  );
  nor  g661( wr_652  , wr_651  , wr_648  );
  not  g662( G72     ,           wr_672  );
  nor  g663( wr_679  , wr_678  , wr_676  );
  nor  g664( wr_589  , wr_588  , G953    );
  nor  g665( wr_603  , wr_602  , wr_599  );
  nor  g666( wr_612  , wr_611  , wr_608  );
  nor  g667( wr_620  , wr_619  , wr_616  );
  nor  g668( wr_628  , wr_627  , wr_624  );
  nor  g669( wr_636  , wr_635  , wr_632  );
  not  g670( G69     ,           wr_652  );
  not  g671( wr_681  ,           wr_679  );
  not  g672( wr_590  ,           wr_589  );
  nor  g673( wr_680  , wr_679  , wr_196  );
  nor  g674( G51     , wr_604  , wr_603  );
  nor  g675( G54     , wr_612  , wr_604  );
  nor  g676( G60     , wr_620  , wr_604  );
  nor  g677( G63     , wr_628  , wr_604  );
  nor  g678( G66     , wr_636  , wr_604  );
  nor  g679( wr_682  , wr_681  , wr_195  );
  nor  g680( wr_591  , wr_590  , wr_492  );
  nor  g681( wr_683  , wr_682  , wr_680  );
  nor  g682( G75     , wr_591  , wr_495  );
  nor  g683( G57     , wr_683  , wr_604  );

endmodule
