// Benchmark "./input/c5315" written by ABC on Thu Aug  8 02:45:58 2024

module c5315  ( 
    G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37,
    G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79,
    G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106,
    G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140,
    G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173,
    G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209,
    G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251,
    G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293,
    G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338,
    G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389,
    G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523,
    G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691,
    G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717,
    G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115,
    G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612,
    G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921,
    G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636,
    G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626,
    G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623,
    G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000,
    G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802,
    G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826,
    G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742,
    G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843,
    G882, G767, G807, G658, G690  );
  input  G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34,
    G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76,
    G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103,
    G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121,
    G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137,
    G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170,
    G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206,
    G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248,
    G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292,
    G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335,
    G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386,
    G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514,
    G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690,
    G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552,
    G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115;
  output G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611,
    G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923,
    G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593,
    G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615,
    G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861,
    G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998,
    G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792,
    G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813,
    G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732,
    G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685,
    G688, G843, G882, G767, G807, G658, G690;
  wire new_G4114_, new_G2825_, new_G3547_, new_G3549_, new_G3551_,
    new_G3553_, new_G633_, new_G814_, new_G816_, new_G844_, new_G846_,
    new_G852_, new_G1502_, new_G1528_, new_G1552_, new_G1609_, new_G1633_,
    new_G1697_, new_G1698_, new_G1701_, new_G2179_, new_G2203_, new_G2226_,
    new_G2281_, new_G2304_, new_G2361_, new_G2370_, new_G2382_, new_G2393_,
    new_G2405_, new_G2418_, new_G2442_, new_G2476_, new_G2500_, new_G2533_,
    new_G2537_, new_G2541_, new_G2545_, new_G2549_, new_G2553_, new_G2557_,
    new_G2561_, new_G2627_, new_G2631_, new_G2635_, new_G2639_, new_G2643_,
    new_G2647_, new_G2651_, new_G2655_, new_G2721_, new_G2734_, new_G2816_,
    new_G2822_, new_G2826_, new_G2828_, new_G2882_, new_G2886_, new_G2890_,
    new_G2894_, new_G2898_, new_G2902_, new_G2948_, new_G2952_, new_G2956_,
    new_G2960_, new_G2964_, new_G2968_, new_G3024_, new_G3028_, new_G3032_,
    new_G3036_, new_G3040_, new_G3044_, new_G3048_, new_G3052_, new_G3092_,
    new_G3105_, new_G3175_, new_G3176_, new_G3181_, new_G3204_, new_G3208_,
    new_G3212_, new_G3216_, new_G3220_, new_G3224_, new_G3256_, new_G3260_,
    new_G3264_, new_G3268_, new_G3272_, new_G3276_, new_G3302_, new_G3314_,
    new_G3354_, new_G3358_, new_G3362_, new_G3366_, new_G3370_, new_G3374_,
    new_G3378_, new_G3382_, new_G3440_, new_G3554_, new_G3555_, new_G3556_,
    new_G3558_, new_G3582_, new_G3616_, new_G3628_, new_G3660_, new_G3684_,
    new_G3721_, new_G3728_, new_G3737_, new_G3757_, new_G3795_, new_G3815_,
    new_G3972_, new_G3991_, new_G4030_, new_G4049_, new_G4110_, new_G4119_,
    new_G4127_, new_G4135_, new_G4143_, new_G4151_, new_G4159_, new_G4167_,
    new_G4175_, new_G4183_, new_G4188_, new_G4276_, new_G4284_, new_G4292_,
    new_G4300_, new_G4308_, new_G4316_, new_G4324_, new_G4332_, new_G4340_,
    new_G4631_, new_G4639_, new_G4647_, new_G4655_, new_G4663_, new_G4671_,
    new_G4676_, new_G4764_, new_G4772_, new_G4780_, new_G4788_, new_G4796_,
    new_G4804_, new_G5082_, new_G5085_, new_G5090_, new_G5093_, new_G5098_,
    new_G5101_, new_G5108_, new_G5111_, new_G5332_, new_G5335_, new_G5340_,
    new_G5343_, new_G5348_, new_G5351_, new_G5356_, new_G5359_, new_G5369_,
    new_G2979_, new_G2999_, new_G1580_, new_G1586_, new_G1592_, new_G1598_,
    new_G1604_, new_G1668_, new_G1674_, new_G1680_, new_G1686_, new_G2254_,
    new_G2260_, new_G2266_, new_G2272_, new_G2278_, new_G2339_, new_G2345_,
    new_G2351_, new_G2357_, new_G711_, new_G721_, new_G726_, new_G731_,
    new_G736_, new_G741_, new_G746_, new_G751_, new_G756_, new_G761_,
    new_G766_, new_G771_, new_G776_, new_G781_, new_G786_, new_G791_,
    new_G796_, new_G801_, new_G806_, new_G3734_, new_G842_, new_G858_,
    new_G881_, new_G4123_, new_G4131_, new_G4139_, new_G4147_, new_G4155_,
    new_G4163_, new_G4171_, new_G4179_, new_G4187_, new_G4194_, new_G4282_,
    new_G4290_, new_G4298_, new_G4306_, new_G4314_, new_G4322_, new_G4330_,
    new_G4338_, new_G4346_, new_G1526_, new_G1540_, new_G1564_, new_G1606_,
    new_G1621_, new_G1645_, new_G1661_, new_G1688_, new_G4635_, new_G4643_,
    new_G4651_, new_G4659_, new_G4667_, new_G4675_, new_G4682_, new_G4770_,
    new_G4778_, new_G4786_, new_G4794_, new_G4802_, new_G4810_, new_G2202_,
    new_G2215_, new_G2238_, new_G2279_, new_G2293_, new_G2316_, new_G2332_,
    new_G2430_, new_G2454_, new_G2488_, new_G2512_, new_G2536_, new_G2540_,
    new_G2544_, new_G2548_, new_G2552_, new_G2556_, new_G2560_, new_G2564_,
    new_G2566_, new_G2572_, new_G2578_, new_G2584_, new_G2590_, new_G2595_,
    new_G2600_, new_G2605_, new_G2630_, new_G2634_, new_G2638_, new_G2642_,
    new_G2646_, new_G2650_, new_G2654_, new_G2658_, new_G2660_, new_G2666_,
    new_G2672_, new_G2678_, new_G2684_, new_G2689_, new_G2694_, new_G2699_,
    new_G2728_, new_G2741_, new_G2748_, new_G2750_, new_G2752_, new_G2754_,
    new_G2756_, new_G2758_, new_G2760_, new_G2762_, new_G2764_, new_G2766_,
    new_G2827_, new_G2838_, new_G2847_, new_G2885_, new_G2889_, new_G2893_,
    new_G2897_, new_G2901_, new_G2905_, new_G2906_, new_G2909_, new_G2913_,
    new_G2918_, new_G2922_, new_G2927_, new_G2951_, new_G2955_, new_G2959_,
    new_G2963_, new_G2967_, new_G2971_, new_G2973_, new_G2980_, new_G2982_,
    new_G2988_, new_G2994_, new_G3001_, new_G3006_, new_G3027_, new_G3031_,
    new_G3035_, new_G3039_, new_G3043_, new_G3047_, new_G3051_, new_G3055_,
    new_G3056_, new_G3060_, new_G3064_, new_G3068_, new_G3073_, new_G3078_,
    new_G3083_, new_G3088_, new_G3099_, new_G3112_, new_G3119_, new_G3121_,
    new_G3123_, new_G3125_, new_G3126_, new_G3128_, new_G3130_, new_G3132_,
    new_G3134_, new_G3136_, new_G3187_, new_G3193_, new_G3196_, new_G3199_,
    new_G3202_, new_G3207_, new_G3211_, new_G3215_, new_G3219_, new_G3223_,
    new_G3227_, new_G3228_, new_G3232_, new_G3234_, new_G3238_, new_G3243_,
    new_G3247_, new_G3249_, new_G3253_, new_G3259_, new_G3263_, new_G3267_,
    new_G3271_, new_G3275_, new_G3279_, new_G3280_, new_G3283_, new_G3287_,
    new_G3292_, new_G3295_, new_G3299_, new_G3305_, new_G3306_, new_G3310_,
    new_G3317_, new_G3318_, new_G3322_, new_G3326_, new_G3333_, new_G3357_,
    new_G3361_, new_G3365_, new_G3369_, new_G3373_, new_G3377_, new_G3381_,
    new_G3385_, new_G3386_, new_G3390_, new_G3394_, new_G3398_, new_G3403_,
    new_G3408_, new_G3413_, new_G3418_, new_G5088_, new_G5089_, new_G5096_,
    new_G5097_, new_G3489_, new_G3493_, new_G3570_, new_G3594_, new_G3622_,
    new_G3632_, new_G3637_, new_G3640_, new_G3643_, new_G3646_, new_G3672_,
    new_G3696_, new_G3745_, new_G3765_, new_G3803_, new_G3823_, new_G5338_,
    new_G5339_, new_G5346_, new_G5347_, new_G5354_, new_G5355_, new_G3979_,
    new_G3998_, new_G4037_, new_G4056_, new_G4094_, new_G5104_, new_G5105_,
    new_G5114_, new_G5115_, new_G5362_, new_G5363_, new_G5366_, new_G5373_,
    new_G2568_, new_G2574_, new_G2580_, new_G2586_, new_G2592_, new_G2597_,
    new_G2602_, new_G2607_, new_G2662_, new_G2668_, new_G2674_, new_G2680_,
    new_G2686_, new_G2691_, new_G2696_, new_G2701_, new_G2907_, new_G2910_,
    new_G2914_, new_G2920_, new_G2924_, new_G2929_, new_G2975_, new_G2984_,
    new_G2990_, new_G2996_, new_G3003_, new_G3008_, new_G3015_, new_G3057_,
    new_G3061_, new_G3065_, new_G3069_, new_G3075_, new_G3080_, new_G3085_,
    new_G3090_, new_G3229_, new_G3233_, new_G3235_, new_G3239_, new_G3244_,
    new_G3250_, new_G3254_, new_G3281_, new_G3284_, new_G3288_, new_G3293_,
    new_G3296_, new_G3300_, new_G3327_, new_G3334_, new_G3387_, new_G3391_,
    new_G3395_, new_G3399_, new_G3405_, new_G3410_, new_G3415_, new_G3420_,
    new_G3422_, new_G3423_, new_G3431_, new_G3432_, new_G3895_, new_G3896_,
    new_G3904_, new_G3905_, new_G3913_, new_G3914_, new_G5106_, new_G5107_,
    new_G5116_, new_G5117_, new_G5364_, new_G5365_, new_G2880_, new_G2881_,
    new_G1579_, new_G1585_, new_G1591_, new_G1597_, new_G1603_, new_G1667_,
    new_G1673_, new_G1679_, new_G1685_, new_G2876_, new_G2877_, new_G2253_,
    new_G2259_, new_G2265_, new_G2271_, new_G2277_, new_G2338_, new_G2344_,
    new_G2350_, new_G2356_, new_G2868_, new_G2869_, new_G710_, new_G2872_,
    new_G2873_, new_G720_, new_G725_, new_G730_, new_G735_, new_G740_,
    new_G745_, new_G750_, new_G755_, new_G760_, new_G765_, new_G770_,
    new_G775_, new_G780_, new_G785_, new_G790_, new_G795_, new_G800_,
    new_G805_, new_G841_, new_G857_, new_G880_, new_G1660_, new_G2331_,
    new_G2569_, new_G2575_, new_G2581_, new_G2587_, new_G2593_, new_G2598_,
    new_G2603_, new_G2608_, new_G2663_, new_G2669_, new_G2675_, new_G2681_,
    new_G2687_, new_G2692_, new_G2697_, new_G2702_, new_G2747_, new_G2749_,
    new_G2751_, new_G2753_, new_G2755_, new_G2757_, new_G2759_, new_G2761_,
    new_G2763_, new_G2765_, new_G2857_, new_G2908_, new_G2911_, new_G2915_,
    new_G2925_, new_G2930_, new_G2933_, new_G2976_, new_G2985_, new_G2991_,
    new_G2997_, new_G3004_, new_G3009_, new_G3058_, new_G3062_, new_G3066_,
    new_G3070_, new_G3076_, new_G3081_, new_G3086_, new_G3091_, new_G3118_,
    new_G3120_, new_G3122_, new_G3124_, new_G3127_, new_G3129_, new_G3131_,
    new_G3133_, new_G3135_, new_G3147_, new_G3192_, new_G3195_, new_G3198_,
    new_G3201_, new_G3230_, new_G3236_, new_G3240_, new_G3245_, new_G3251_,
    new_G3255_, new_G3282_, new_G3285_, new_G3289_, new_G3297_, new_G3301_,
    new_G3309_, new_G3313_, new_G3321_, new_G3325_, new_G3328_, new_G3329_,
    new_G3335_, new_G3336_, new_G3341_, new_G3345_, new_G3388_, new_G3392_,
    new_G3396_, new_G3400_, new_G3406_, new_G3411_, new_G3416_, new_G3421_,
    new_G3424_, new_G3433_, new_G3492_, new_G3496_, new_G3780_, new_G3783_,
    new_G3786_, new_G3789_, new_G3838_, new_G3841_, new_G3844_, new_G3847_,
    new_G3897_, new_G3906_, new_G3915_, new_G4011_, new_G4014_, new_G4017_,
    new_G4020_, new_G4023_, new_G4069_, new_G4072_, new_G4075_, new_G4078_,
    new_G4081_, new_G5206_, new_G5209_, new_G5307_, new_G5322_, new_G5372_,
    new_G5375_, new_G5399_, new_G2813_, new_G3197_, new_G3200_, new_G3203_,
    new_G3194_, new_G2570_, new_G2576_, new_G2582_, new_G2588_, new_G2664_,
    new_G2670_, new_G2676_, new_G2682_, new_G2767_, new_G2772_, new_G2776_,
    new_G2780_, new_G2784_, new_G2788_, new_G2794_, new_G2798_, new_G2802_,
    new_G2912_, new_G2916_, new_G2936_, new_G2977_, new_G2986_, new_G2992_,
    new_G3059_, new_G3063_, new_G3067_, new_G3071_, new_G3137_, new_G3139_,
    new_G3143_, new_G3151_, new_G3155_, new_G3161_, new_G3165_, new_G3167_,
    new_G3231_, new_G3237_, new_G3241_, new_G3286_, new_G3290_, new_G3330_,
    new_G3337_, new_G3342_, new_G3346_, new_G3348_, new_G3352_, new_G3389_,
    new_G3393_, new_G3397_, new_G3401_, new_G3845_, new_G5126_, new_G5178_,
    new_G5325_, new_G5374_, new_G2810_, new_G635_, new_G2878_, new_G2879_,
    new_G2874_, new_G2875_, new_G703_, new_G2866_, new_G2867_, new_G2870_,
    new_G2871_, new_G716_, new_G819_, new_G1789_, new_G2036_, new_G2611_,
    new_G2615_, new_G2619_, new_G2623_, new_G2705_, new_G2709_, new_G2713_,
    new_G2717_, new_G2939_, new_G2942_, new_G2945_, new_G3012_, new_G3018_,
    new_G3021_, new_G3331_, new_G3338_, new_G3343_, new_G3347_, new_G3428_,
    new_G3437_, new_G3514_, new_G3836_, new_G3852_, new_G5311_, new_G3901_,
    new_G3910_, new_G3934_, new_G3938_, new_G4652_, new_G4783_, new_G5137_,
    new_G5212_, new_G5213_, new_G5260_, new_G5263_, new_G5268_, new_G5271_,
    new_G5276_, new_G5279_, new_G5289_, new_G5296_, new_G5299_, new_G5304_,
    new_G5312_, new_G5315_, new_G5328_, new_G5396_, new_G5403_, new_G1286_,
    new_G2809_, new_G597_, new_G1031_, new_G637_, new_G671_, new_G705_,
    new_G713_, new_G1046_, new_G1064_, new_G1071_, new_G1097_, new_G1111_,
    new_G1128_, new_G1145_, new_G1160_, new_G1301_, new_G1318_, new_G1324_,
    new_G1341_, new_G1359_, new_G1382_, new_G1404_, new_G1412_, new_G1704_,
    new_G1712_, new_G1724_, new_G1742_, new_G1749_, new_G1775_, new_G1806_,
    new_G1823_, new_G1829_, new_G1837_, new_G1958_, new_G1966_, new_G1978_,
    new_G1995_, new_G2001_, new_G2018_, new_G2059_, new_G2081_, new_G2089_,
    new_G2106_, new_G3170_, new_G3332_, new_G3339_, new_G5132_, new_G5184_,
    new_G3853_, new_G3874_, new_G4076_, new_G4116_, new_G4124_, new_G4132_,
    new_G4140_, new_G4148_, new_G4156_, new_G4164_, new_G4172_, new_G4180_,
    new_G4228_, new_G4279_, new_G4287_, new_G4295_, new_G4303_, new_G4311_,
    new_G4319_, new_G4327_, new_G4335_, new_G4343_, new_G4348_, new_G4464_,
    new_G4628_, new_G4636_, new_G4644_, new_G4660_, new_G4668_, new_G4716_,
    new_G4767_, new_G4775_, new_G4791_, new_G4799_, new_G4807_, new_G4812_,
    new_G5118_, new_G5121_, new_G5129_, new_G5134_, new_G5142_, new_G5145_,
    new_G5152_, new_G5155_, new_G5162_, new_G5165_, new_G5170_, new_G5173_,
    new_G5181_, new_G5186_, new_G5189_, new_G5196_, new_G5199_, new_G5214_,
    new_G5215_, new_G5329_, new_G5330_, new_G2807_, new_G2808_, new_G2811_,
    new_G2812_, new_G2814_, new_G2626_, new_G2622_, new_G2618_, new_G2614_,
    new_G2720_, new_G2716_, new_G2712_, new_G2708_, new_G3731_, new_G4658_,
    new_G1777_, new_G2019_, new_G4787_, new_G3350_, new_G3353_, new_G5141_,
    new_G3513_, new_G3516_, new_G3517_, new_G3778_, new_G3781_, new_G3784_,
    new_G3787_, new_G3839_, new_G3842_, new_G5266_, new_G5267_, new_G5274_,
    new_G5275_, new_G5302_, new_G5303_, new_G5310_, new_G3891_, new_G3937_,
    new_G3941_, new_G3955_, new_G3958_, new_G4009_, new_G4012_, new_G4015_,
    new_G4018_, new_G4067_, new_G4070_, new_G4073_, new_G4079_, new_G5239_,
    new_G5282_, new_G5283_, new_G5293_, new_G5318_, new_G5319_, new_G5331_,
    new_G5402_, new_G5405_, new_G595_, new_G596_, new_G607_, new_G608_,
    new_G1845_, new_G1846_, new_G2115_, new_G2116_, new_G4122_, new_G1022_,
    new_G4130_, new_G1033_, new_G4138_, new_G1051_, new_G4146_, new_G1079_,
    new_G4154_, new_G1088_, new_G4162_, new_G1099_, new_G4170_, new_G1115_,
    new_G4178_, new_G1133_, new_G4186_, new_G1151_, new_G4234_, new_G1276_,
    new_G4283_, new_G1287_, new_G4291_, new_G1305_, new_G4299_, new_G1330_,
    new_G4307_, new_G1342_, new_G4315_, new_G1363_, new_G4323_, new_G1388_,
    new_G4331_, new_G1420_, new_G4339_, new_G1428_, new_G4347_, new_G4634_,
    new_G1729_, new_G4642_, new_G1757_, new_G4650_, new_G1766_, new_G1776_,
    new_G4666_, new_G1793_, new_G4674_, new_G1811_, new_G1849_, new_G1852_,
    new_G1875_, new_G4722_, new_G1982_, new_G4771_, new_G2007_, new_G4779_,
    new_G2020_, new_G2040_, new_G4795_, new_G2065_, new_G4803_, new_G2097_,
    new_G4811_, new_G2119_, new_G2122_, new_G5124_, new_G5125_, new_G3452_,
    new_G5133_, new_G5140_, new_G3462_, new_G5168_, new_G5169_, new_G5176_,
    new_G5177_, new_G3484_, new_G5185_, new_G3515_, new_G3518_, new_G3857_,
    new_G3860_, new_G3861_, new_G3869_, new_G3870_, new_G3878_, new_G3881_,
    new_G3882_, new_G3890_, new_G3954_, new_G3957_, new_G4021_, new_G4099_,
    new_G4236_, new_G4354_, new_G4406_, new_G4470_, new_G4552_, new_G4679_,
    new_G4687_, new_G4695_, new_G4703_, new_G4711_, new_G4724_, new_G4818_,
    new_G4855_, new_G4865_, new_G4870_, new_G4913_, new_G4923_, new_G4951_,
    new_G5006_, new_G5039_, new_G5148_, new_G5149_, new_G5158_, new_G5159_,
    new_G5192_, new_G5193_, new_G5202_, new_G5203_, new_G5284_, new_G5285_,
    new_G5320_, new_G5321_, new_G5386_, new_G5404_, new_G609_, new_G1021_,
    new_G1032_, new_G1050_, new_G1078_, new_G1087_, new_G1098_, new_G1114_,
    new_G1132_, new_G1150_, new_G1277_, new_G1288_, new_G1306_, new_G1331_,
    new_G1343_, new_G1364_, new_G1389_, new_G1421_, new_G1429_, new_G1728_,
    new_G1756_, new_G1765_, new_G1778_, new_G1792_, new_G1810_, new_G1983_,
    new_G2008_, new_G2021_, new_G2041_, new_G2066_, new_G2098_, new_G3443_,
    new_G3444_, new_G3453_, new_G3461_, new_G3466_, new_G3467_, new_G3475_,
    new_G3476_, new_G3485_, new_G5243_, new_G3862_, new_G3871_, new_G3883_,
    new_G3892_, new_G3956_, new_G3959_, new_G4756_, new_G5150_, new_G5151_,
    new_G5160_, new_G5161_, new_G5194_, new_G5195_, new_G5204_, new_G5205_,
    new_G5236_, new_G5286_, new_G5379_, new_G5389_, new_G5425_, new_G1023_,
    new_G1034_, new_G1052_, new_G1080_, new_G1089_, new_G1100_, new_G1116_,
    new_G1134_, new_G1152_, new_G4242_, new_G1278_, new_G1289_, new_G1307_,
    new_G1332_, new_G1344_, new_G1365_, new_G1390_, new_G1422_, new_G1430_,
    new_G1730_, new_G1758_, new_G1767_, new_G1794_, new_G1812_, new_G1876_,
    new_G4683_, new_G4691_, new_G4699_, new_G4707_, new_G4715_, new_G4730_,
    new_G1984_, new_G2009_, new_G2042_, new_G2067_, new_G2099_, new_G4869_,
    new_G4927_, new_G3445_, new_G3454_, new_G3463_, new_G3468_, new_G3477_,
    new_G3486_, new_G4103_, new_G4412_, new_G4558_, new_G4859_, new_G4876_,
    new_G4917_, new_G4955_, new_G5012_, new_G5043_, new_G5216_, new_G5219_,
    new_G5226_, new_G5229_, new_G5392_, new_G5422_, new_G1866_, new_G1877_,
    new_G4762_, new_G2142_, new_G2146_, new_G5242_, new_G3532_, new_G3866_,
    new_G3887_, new_G3918_, new_G3922_, new_G3926_, new_G3930_, new_G5429_,
    new_G4104_, new_G4743_, new_G4991_, new_G5001_, new_G5292_, new_G5295_,
    new_G5383_, new_G5393_, new_G5394_, new_G1439_, new_G1440_, new_G1441_,
    new_G1847_, new_G1168_, new_G1169_, new_G1170_, new_G2117_, new_G1086_,
    new_G1166_, new_G1171_, new_G1172_, new_G1173_, new_G1174_, new_G1175_,
    new_G1176_, new_G1177_, new_G1178_, new_G1179_, new_G1181_, new_G1182_,
    new_G1183_, new_G1184_, new_G1188_, new_G1189_, new_G1190_, new_G1191_,
    new_G1192_, new_G1193_, new_G1194_, new_G1195_, new_G1196_, new_G1197_,
    new_G1437_, new_G1442_, new_G1443_, new_G1444_, new_G1445_, new_G1446_,
    new_G1447_, new_G1451_, new_G1454_, new_G1455_, new_G1456_, new_G1457_,
    new_G1465_, new_G1466_, new_G1467_, new_G1468_, new_G1469_, new_G1470_,
    new_G1471_, new_G1472_, new_G1473_, new_G1474_, new_G1475_, new_G1476_,
    new_G1477_, new_G1481_, new_G1482_, new_G1764_, new_G1843_, new_G1850_,
    new_G1851_, new_G1853_, new_G1854_, new_G1855_, new_G1856_, new_G1857_,
    new_G1859_, new_G1860_, new_G1861_, new_G1862_, new_G1867_, new_G1868_,
    new_G1869_, new_G1870_, new_G1871_, new_G1872_, new_G1873_, new_G1874_,
    new_G1878_, new_G2113_, new_G2120_, new_G2121_, new_G2123_, new_G2124_,
    new_G2128_, new_G2131_, new_G2132_, new_G2133_, new_G2134_, new_G2143_,
    new_G2144_, new_G2145_, new_G2147_, new_G2148_, new_G2149_, new_G2150_,
    new_G2151_, new_G2152_, new_G2153_, new_G2154_, new_G2158_, new_G2159_,
    new_G3449_, new_G3458_, new_G3472_, new_G3481_, new_G3497_, new_G3501_,
    new_G3505_, new_G3509_, new_G3531_, new_G5428_, new_G3967_, new_G4191_,
    new_G4199_, new_G4207_, new_G4215_, new_G4223_, new_G4231_, new_G4239_,
    new_G4247_, new_G4255_, new_G4263_, new_G4271_, new_G4371_, new_G4381_,
    new_G4391_, new_G4401_, new_G4429_, new_G4439_, new_G4449_, new_G4459_,
    new_G4497_, new_G4507_, new_G4517_, new_G4527_, new_G4537_, new_G4547_,
    new_G4585_, new_G4595_, new_G4605_, new_G4615_, new_G4719_, new_G4727_,
    new_G4735_, new_G4751_, new_G4759_, new_G4835_, new_G4845_, new_G4893_,
    new_G4903_, new_G4961_, new_G4971_, new_G4981_, new_G5049_, new_G5059_,
    new_G5069_, new_G5222_, new_G5223_, new_G5232_, new_G5233_, new_G5294_,
    new_G5395_, new_G589_, new_G616_, new_G619_, new_G627_, new_G1185_,
    new_G1448_, new_G1458_, new_G1478_, new_G1863_, new_G4747_, new_G2125_,
    new_G2135_, new_G2155_, new_G4995_, new_G5005_, new_G3533_, new_G3921_,
    new_G3925_, new_G3929_, new_G3933_, new_G3943_, new_G3946_, new_G3949_,
    new_G3952_, new_G3966_, new_G4107_, new_G4196_, new_G4204_, new_G4212_,
    new_G4220_, new_G4244_, new_G4252_, new_G4260_, new_G4268_, new_G4361_,
    new_G4419_, new_G4467_, new_G4487_, new_G4555_, new_G4575_, new_G4684_,
    new_G4692_, new_G4700_, new_G4708_, new_G4732_, new_G4740_, new_G4748_,
    new_G4825_, new_G4883_, new_G4928_, new_G4941_, new_G5009_, new_G5029_,
    new_G5224_, new_G5225_, new_G5234_, new_G5235_, new_G5376_, new_G5417_,
    new_G576_, new_G1198_, new_G4195_, new_G4203_, new_G4211_, new_G4219_,
    new_G4227_, new_G1217_, new_G4235_, new_G1221_, new_G4243_, new_G1224_,
    new_G4251_, new_G4259_, new_G4267_, new_G4275_, new_G1453_, new_G4405_,
    new_G4463_, new_G4541_, new_G4551_, new_G1895_, new_G4723_, new_G1899_,
    new_G4731_, new_G1902_, new_G4739_, new_G4755_, new_G1929_, new_G4763_,
    new_G2130_, new_G3500_, new_G3504_, new_G3508_, new_G3512_, new_G3520_,
    new_G3523_, new_G3526_, new_G3529_, new_G3837_, new_G3942_, new_G3945_,
    new_G3948_, new_G3951_, new_G3968_, new_G4375_, new_G4385_, new_G4395_,
    new_G4433_, new_G4443_, new_G4453_, new_G4501_, new_G4511_, new_G4521_,
    new_G4531_, new_G4619_, new_G4589_, new_G4599_, new_G4609_, new_G4839_,
    new_G4849_, new_G4897_, new_G4907_, new_G4965_, new_G4975_, new_G4985_,
    new_G5073_, new_G5053_, new_G5063_, new_G5247_, new_G5255_, new_G590_,
    new_G617_, new_G620_, new_G628_, new_G3535_, new_G1199_, new_G4202_,
    new_G1204_, new_G4210_, new_G1207_, new_G4218_, new_G1211_, new_G4226_,
    new_G1214_, new_G1218_, new_G1222_, new_G1225_, new_G4250_, new_G1237_,
    new_G4258_, new_G1242_, new_G4266_, new_G1247_, new_G4274_, new_G1252_,
    new_G1462_, new_G4690_, new_G1882_, new_G4698_, new_G1885_, new_G4706_,
    new_G1889_, new_G4714_, new_G1892_, new_G1896_, new_G1900_, new_G1903_,
    new_G4738_, new_G1915_, new_G4746_, new_G1920_, new_G4754_, new_G1925_,
    new_G1930_, new_G2139_, new_G3519_, new_G3522_, new_G3525_, new_G3528_,
    new_G3848_, new_G3944_, new_G3947_, new_G3950_, new_G3953_, new_G5421_,
    new_G4111_, new_G4112_, new_G4351_, new_G4365_, new_G4409_, new_G4423_,
    new_G4471_, new_G4472_, new_G4477_, new_G4491_, new_G4559_, new_G4560_,
    new_G4565_, new_G4579_, new_G4815_, new_G4829_, new_G4873_, new_G4887_,
    new_G4931_, new_G4934_, new_G4945_, new_G5013_, new_G5014_, new_G5019_,
    new_G5033_, new_G5382_, new_G5385_, new_G3970_, new_G1200_, new_G1203_,
    new_G1206_, new_G1210_, new_G1213_, new_G1219_, new_G1223_, new_G1236_,
    new_G1241_, new_G1246_, new_G1251_, new_G1881_, new_G1884_, new_G1888_,
    new_G1891_, new_G1897_, new_G1901_, new_G1914_, new_G1919_, new_G1924_,
    new_G1931_, new_G3521_, new_G3524_, new_G3527_, new_G3530_, new_G5251_,
    new_G5259_, new_G4113_, new_G4473_, new_G4561_, new_G5015_, new_G5384_,
    new_G5406_, new_G5414_, new_G1664_, new_G2335_, new_G718_, new_G855_,
    new_G1205_, new_G1208_, new_G1212_, new_G1215_, new_G1220_, new_G1231_,
    new_G1238_, new_G1243_, new_G1248_, new_G1253_, new_G1272_, new_G1483_,
    new_G1883_, new_G1886_, new_G1890_, new_G1893_, new_G1898_, new_G1909_,
    new_G1916_, new_G1921_, new_G1926_, new_G1953_, new_G2160_, new_G4355_,
    new_G4356_, new_G4413_, new_G4414_, new_G4474_, new_G4481_, new_G4562_,
    new_G4569_, new_G4819_, new_G4820_, new_G4877_, new_G4878_, new_G4935_,
    new_G4936_, new_G5016_, new_G5023_, new_G5244_, new_G5252_, new_G5409_,
    new_G566_, new_G577_, new_G3733_, new_G1209_, new_G1216_, new_G1257_,
    new_G1262_, new_G1267_, new_G1887_, new_G1894_, new_G1935_, new_G1943_,
    new_G1948_, new_G3779_, new_G3840_, new_G5412_, new_G5420_, new_G3964_,
    new_G4357_, new_G4415_, new_G4821_, new_G4879_, new_G4937_, new_G567_,
    new_G568_, new_G569_, new_G570_, new_G578_, new_G579_, new_G580_,
    new_G1256_, new_G1261_, new_G1266_, new_G1271_, new_G1486_, new_G1934_,
    new_G1942_, new_G1947_, new_G1952_, new_G2163_, new_G5250_, new_G3537_,
    new_G5258_, new_G3542_, new_G3782_, new_G3785_, new_G3788_, new_G3790_,
    new_G3843_, new_G3846_, new_G3849_, new_G3960_, new_G5413_, new_G3963_,
    new_G4010_, new_G4068_, new_G4358_, new_G4416_, new_G4480_, new_G4483_,
    new_G4568_, new_G4571_, new_G4822_, new_G4880_, new_G4938_, new_G5022_,
    new_G5025_, new_G1258_, new_G1263_, new_G1268_, new_G1273_, new_G1936_,
    new_G1944_, new_G1949_, new_G1954_, new_G3536_, new_G3541_, new_G3791_,
    new_G3792_, new_G3793_, new_G3850_, new_G3851_, new_G3961_, new_G3965_,
    new_G4024_, new_G4082_, new_G4482_, new_G4570_, new_G5024_, new_G1666_,
    new_G1670_, new_G2337_, new_G2341_, new_G719_, new_G758_, new_G798_,
    new_G856_, new_G3538_, new_G3543_, new_G3962_, new_G4364_, new_G4367_,
    new_G4422_, new_G4425_, new_G4484_, new_G4572_, new_G4828_, new_G4831_,
    new_G4886_, new_G4889_, new_G4944_, new_G4947_, new_G5026_, new_G571_,
    new_G572_, new_G573_, new_G574_, new_G581_, new_G582_, new_G583_,
    new_G584_, new_G1576_, new_G1578_, new_G659_, new_G1672_, new_G1676_,
    new_G1678_, new_G1682_, new_G1684_, new_G2250_, new_G2252_, new_G691_,
    new_G2343_, new_G2347_, new_G2349_, new_G2353_, new_G2355_, new_G743_,
    new_G744_, new_G748_, new_G749_, new_G753_, new_G754_, new_G759_,
    new_G783_, new_G784_, new_G788_, new_G789_, new_G793_, new_G794_,
    new_G799_, new_G3735_, new_G3835_, new_G3651_, new_G4013_, new_G4016_,
    new_G4019_, new_G4022_, new_G4071_, new_G4074_, new_G4077_, new_G4080_,
    new_G4096_, new_G4366_, new_G4424_, new_G4830_, new_G4888_, new_G4946_,
    new_G640_, new_G662_, new_G665_, new_G668_, new_G674_, new_G694_,
    new_G697_, new_G700_, new_G817_, new_G839_, new_G3540_, new_G3545_,
    new_G3777_, new_G3648_, new_G4025_, new_G4026_, new_G4027_, new_G4028_,
    new_G4083_, new_G4084_, new_G4085_, new_G4086_, new_G4368_, new_G4426_,
    new_G4490_, new_G4493_, new_G4578_, new_G4581_, new_G4832_, new_G4890_,
    new_G4948_, new_G5032_, new_G5035_, new_G811_, new_G812_, new_G853_,
    new_G878_, new_G4492_, new_G4580_, new_G5034_, new_G1582_, new_G1584_,
    new_G1588_, new_G1590_, new_G1594_, new_G1596_, new_G1600_, new_G1602_,
    new_G2256_, new_G2258_, new_G2262_, new_G2264_, new_G2268_, new_G2270_,
    new_G2274_, new_G2276_, new_G708_, new_G709_, new_G723_, new_G724_,
    new_G728_, new_G729_, new_G733_, new_G734_, new_G738_, new_G739_,
    new_G768_, new_G769_, new_G773_, new_G774_, new_G778_, new_G779_,
    new_G4374_, new_G4377_, new_G4432_, new_G4435_, new_G4494_, new_G4582_,
    new_G4838_, new_G4841_, new_G4896_, new_G4899_, new_G4954_, new_G4957_,
    new_G5036_, new_G643_, new_G646_, new_G649_, new_G652_, new_G677_,
    new_G680_, new_G683_, new_G686_, new_G4376_, new_G4434_, new_G4840_,
    new_G4898_, new_G4956_, new_G4378_, new_G4436_, new_G4500_, new_G4503_,
    new_G4588_, new_G4591_, new_G4842_, new_G4900_, new_G4958_, new_G5042_,
    new_G5045_, new_G4502_, new_G4590_, new_G5044_, new_G4384_, new_G4387_,
    new_G4442_, new_G4445_, new_G4504_, new_G4592_, new_G4848_, new_G4851_,
    new_G4906_, new_G4909_, new_G4964_, new_G4967_, new_G5046_, new_G4386_,
    new_G4444_, new_G4850_, new_G4908_, new_G4966_, new_G4388_, new_G4446_,
    new_G4510_, new_G4513_, new_G4598_, new_G4601_, new_G4852_, new_G4910_,
    new_G4968_, new_G5052_, new_G5055_, new_G4512_, new_G4600_, new_G5054_,
    new_G4394_, new_G4397_, new_G4452_, new_G4455_, new_G4514_, new_G4602_,
    new_G4858_, new_G4861_, new_G4916_, new_G4919_, new_G4974_, new_G4977_,
    new_G5056_, new_G4396_, new_G4454_, new_G4860_, new_G4918_, new_G4976_,
    new_G4398_, new_G4456_, new_G4520_, new_G4523_, new_G4608_, new_G4611_,
    new_G4862_, new_G4920_, new_G4978_, new_G5062_, new_G5065_, new_G4522_,
    new_G4610_, new_G5064_, new_G4404_, new_G1488_, new_G4462_, new_G1493_,
    new_G4868_, new_G2165_, new_G4926_, new_G2170_, new_G4524_, new_G4612_,
    new_G4984_, new_G4987_, new_G5066_, new_G1487_, new_G1492_, new_G2164_,
    new_G2169_, new_G4986_, new_G1489_, new_G1494_, new_G2166_, new_G2171_,
    new_G4530_, new_G4533_, new_G4618_, new_G4543_, new_G4988_, new_G5072_,
    new_G4997_, new_G4532_, new_G4542_, new_G4996_, new_G1513_, new_G1514_,
    new_G1515_, new_G1516_, new_G4994_, new_G2184_, new_G2190_, new_G2191_,
    new_G2192_, new_G2193_, new_G4534_, new_G4544_, new_G4998_, new_G2183_,
    new_G4620_, new_G5074_, new_G4540_, new_G1507_, new_G4550_, new_G1510_,
    new_G2185_, new_G5004_, new_G2187_, new_G1506_, new_G1509_, new_G4626_,
    new_G2186_, new_G2195_, new_G5080_, new_G1508_, new_G1511_, new_G2188_,
    new_G1512_, new_G1518_, new_G2189_, new_G1517_, new_G2194_, new_G4623_,
    new_G5077_, new_G1519_, new_G4627_, new_G2196_, new_G5081_, new_G1520_,
    new_G2197_, new_G1521_, new_G2198_, new_G840_, new_G879_, new_G1524_,
    new_G2201_, new_G3649_, new_G3652_, new_G3657_, new_G3658_, new_G3636_,
    new_G3639_, new_G3642_, new_G3645_, new_G3653_, new_G3654_, new_G3655_,
    new_G3656_, new_G763_, new_G764_, new_G803_, new_G804_, new_G1657_,
    new_G1659_, new_G2328_, new_G2330_, new_G1662_, new_G2333_, new_G657_,
    new_G689_;
  assign G144 = G141;
  assign G298 = G293;
  assign new_G4114_ = G135 & G4115;
  assign new_G2825_ = ~G2824;
  assign G973 = G3173;
  assign new_G3547_ = ~G3546;
  assign new_G3549_ = ~G3548;
  assign new_G3551_ = ~G3550;
  assign new_G3553_ = ~G3552;
  assign G594 = ~G545;
  assign G599 = ~G348;
  assign G600 = ~G366;
  assign G601 = G552 & G562;
  assign G602 = ~G549;
  assign G603 = ~G545;
  assign G604 = ~G545;
  assign G611 = ~G338;
  assign G612 = ~G358;
  assign new_G633_ = ~G373 | ~G1;
  assign G810 = G141 & G145;
  assign new_G814_ = ~G3173;
  assign new_G816_ = ~new_G4114_;
  assign new_G844_ = new_G2825_ & G27;
  assign new_G846_ = G386 & G556;
  assign G848 = ~G245;
  assign G849 = ~G552;
  assign G850 = ~G562;
  assign G851 = ~G559;
  assign new_G852_ = G552 & G556 & G386 & G559;
  assign new_G1502_ = ~G1497;
  assign new_G1528_ = G1689;
  assign new_G1552_ = G1690;
  assign new_G1609_ = G1689;
  assign new_G1633_ = G1690;
  assign new_G1697_ = G137;
  assign new_G1698_ = G137;
  assign new_G1701_ = G141;
  assign new_G2179_ = ~G2174;
  assign new_G2203_ = G1691;
  assign new_G2226_ = G1694;
  assign new_G2281_ = G1691;
  assign new_G2304_ = G1694;
  assign new_G2361_ = G254;
  assign new_G2370_ = G251;
  assign new_G2382_ = G251;
  assign new_G2393_ = G248;
  assign new_G2405_ = G248;
  assign new_G2418_ = G4088;
  assign new_G2442_ = G4087;
  assign new_G2476_ = G4089;
  assign new_G2500_ = G4090;
  assign new_G2533_ = G210;
  assign new_G2537_ = G210;
  assign new_G2541_ = G218;
  assign new_G2545_ = G218;
  assign new_G2549_ = G226;
  assign new_G2553_ = G226;
  assign new_G2557_ = G234;
  assign new_G2561_ = G234;
  assign new_G2627_ = G257;
  assign new_G2631_ = G257;
  assign new_G2635_ = G265;
  assign new_G2639_ = G265;
  assign new_G2643_ = G273;
  assign new_G2647_ = G273;
  assign new_G2651_ = G281;
  assign new_G2655_ = G281;
  assign new_G2721_ = G335;
  assign new_G2734_ = G335;
  assign new_G2816_ = G206;
  assign new_G2822_ = G27 & G31;
  assign new_G2826_ = G1;
  assign new_G2828_ = G2358;
  assign new_G2882_ = G293;
  assign new_G2886_ = G302;
  assign new_G2890_ = G308;
  assign new_G2894_ = G308;
  assign new_G2898_ = G316;
  assign new_G2902_ = G316;
  assign new_G2948_ = G324;
  assign new_G2952_ = G324;
  assign new_G2956_ = G341;
  assign new_G2960_ = G341;
  assign new_G2964_ = G351;
  assign new_G2968_ = G351;
  assign new_G3024_ = G257;
  assign new_G3028_ = G257;
  assign new_G3032_ = G265;
  assign new_G3036_ = G265;
  assign new_G3040_ = G273;
  assign new_G3044_ = G273;
  assign new_G3048_ = G281;
  assign new_G3052_ = G281;
  assign new_G3092_ = G332;
  assign new_G3105_ = G332;
  assign new_G3175_ = G549;
  assign new_G3176_ = G31 & G27;
  assign new_G3181_ = ~G2358;
  assign new_G3204_ = G324;
  assign new_G3208_ = G324;
  assign new_G3212_ = G341;
  assign new_G3216_ = G341;
  assign new_G3220_ = G351;
  assign new_G3224_ = G351;
  assign new_G3256_ = G293;
  assign new_G3260_ = G302;
  assign new_G3264_ = G308;
  assign new_G3268_ = G308;
  assign new_G3272_ = G316;
  assign new_G3276_ = G316;
  assign new_G3302_ = G361;
  assign new_G3314_ = G361;
  assign new_G3354_ = G210;
  assign new_G3358_ = G210;
  assign new_G3362_ = G218;
  assign new_G3366_ = G218;
  assign new_G3370_ = G226;
  assign new_G3374_ = G226;
  assign new_G3378_ = G234;
  assign new_G3382_ = G234;
  assign new_G3440_ = ~G324;
  assign new_G3554_ = G242;
  assign new_G3555_ = G242;
  assign new_G3556_ = G254;
  assign new_G3558_ = G4088;
  assign new_G3582_ = G4087;
  assign new_G3616_ = G4092;
  assign new_G3628_ = G4091;
  assign new_G3660_ = G4089;
  assign new_G3684_ = G4090;
  assign new_G3721_ = ~G3717;
  assign new_G3728_ = ~G3724;
  assign new_G3737_ = G4091;
  assign new_G3757_ = G4092;
  assign new_G3795_ = G4091;
  assign new_G3815_ = G4092;
  assign new_G3972_ = G4091;
  assign new_G3991_ = G4092;
  assign new_G4030_ = G4091;
  assign new_G4049_ = G4092;
  assign new_G4110_ = G299;
  assign new_G4119_ = G446;
  assign new_G4127_ = G457;
  assign new_G4135_ = G468;
  assign new_G4143_ = G422;
  assign new_G4151_ = G435;
  assign new_G4159_ = G389;
  assign new_G4167_ = G400;
  assign new_G4175_ = G411;
  assign new_G4183_ = G374;
  assign new_G4188_ = G4;
  assign new_G4276_ = G446;
  assign new_G4284_ = G457;
  assign new_G4292_ = G468;
  assign new_G4300_ = G435;
  assign new_G4308_ = G389;
  assign new_G4316_ = G400;
  assign new_G4324_ = G411;
  assign new_G4332_ = G422;
  assign new_G4340_ = G374;
  assign new_G4631_ = G479;
  assign new_G4639_ = G490;
  assign new_G4647_ = G503;
  assign new_G4655_ = G514;
  assign new_G4663_ = G523;
  assign new_G4671_ = G534;
  assign new_G4676_ = G54;
  assign new_G4764_ = G479;
  assign new_G4772_ = G503;
  assign new_G4780_ = G514;
  assign new_G4788_ = G523;
  assign new_G4796_ = G534;
  assign new_G4804_ = G490;
  assign new_G5082_ = G361;
  assign new_G5085_ = G369;
  assign new_G5090_ = G341;
  assign new_G5093_ = G351;
  assign new_G5098_ = G308;
  assign new_G5101_ = G316;
  assign new_G5108_ = G293;
  assign new_G5111_ = G302;
  assign new_G5332_ = G281;
  assign new_G5335_ = G289;
  assign new_G5340_ = G265;
  assign new_G5343_ = G273;
  assign new_G5348_ = G234;
  assign new_G5351_ = G257;
  assign new_G5356_ = G218;
  assign new_G5359_ = G226;
  assign new_G5369_ = G210;
  assign G634 = ~new_G633_;
  assign G815 = G136 & new_G814_;
  assign G845 = ~new_G844_;
  assign G847 = ~new_G846_;
  assign G926 = new_G1697_;
  assign G923 = new_G1701_;
  assign G921 = new_G2826_;
  assign new_G2979_ = new_G3553_ & G514;
  assign new_G2999_ = new_G3547_ | G514;
  assign G892 = new_G3175_;
  assign G887 = new_G4110_;
  assign G606 = ~new_G3175_;
  assign new_G1580_ = new_G1552_ & G170 & new_G1528_;
  assign new_G1586_ = new_G1552_ & G173 & new_G1528_;
  assign new_G1592_ = new_G1552_ & G167 & new_G1528_;
  assign new_G1598_ = new_G1552_ & G164 & new_G1528_;
  assign new_G1604_ = new_G1552_ & G161 & new_G1528_;
  assign G656 = ~new_G2822_ | ~G140;
  assign new_G1668_ = new_G1633_ & G185 & new_G1609_;
  assign new_G1674_ = new_G1633_ & G158 & new_G1609_;
  assign new_G1680_ = new_G1633_ & G152 & new_G1609_;
  assign new_G1686_ = new_G1633_ & G146 & new_G1609_;
  assign new_G2254_ = new_G2226_ & G170 & new_G2203_;
  assign new_G2260_ = new_G2226_ & G173 & new_G2203_;
  assign new_G2266_ = new_G2226_ & G167 & new_G2203_;
  assign new_G2272_ = new_G2226_ & G164 & new_G2203_;
  assign new_G2278_ = new_G2226_ & G161 & new_G2203_;
  assign new_G2339_ = new_G2304_ & G185 & new_G2281_;
  assign new_G2345_ = new_G2304_ & G158 & new_G2281_;
  assign new_G2351_ = new_G2304_ & G152 & new_G2281_;
  assign new_G2357_ = new_G2304_ & G146 & new_G2281_;
  assign new_G711_ = new_G3684_ & G106 & new_G3660_;
  assign new_G721_ = new_G2442_ & G61 & new_G2418_;
  assign new_G726_ = new_G3582_ & G106 & new_G3558_;
  assign new_G731_ = new_G3582_ & G49 & new_G3558_;
  assign new_G736_ = new_G3582_ & G103 & new_G3558_;
  assign new_G741_ = new_G3582_ & G40 & new_G3558_;
  assign new_G746_ = new_G3582_ & G37 & new_G3558_;
  assign new_G751_ = new_G2442_ & G20 & new_G2418_;
  assign new_G756_ = new_G2442_ & G17 & new_G2418_;
  assign new_G761_ = new_G2442_ & G70 & new_G2418_;
  assign new_G766_ = new_G2442_ & G64 & new_G2418_;
  assign new_G771_ = new_G3684_ & G49 & new_G3660_;
  assign new_G776_ = new_G3684_ & G103 & new_G3660_;
  assign new_G781_ = new_G3684_ & G40 & new_G3660_;
  assign new_G786_ = new_G3684_ & G37 & new_G3660_;
  assign new_G791_ = new_G2500_ & G20 & new_G2476_;
  assign new_G796_ = new_G2500_ & G17 & new_G2476_;
  assign new_G801_ = new_G2500_ & G70 & new_G2476_;
  assign new_G806_ = new_G2500_ & G64 & new_G2476_;
  assign G809 = ~new_G2822_;
  assign new_G3734_ = G3717 & G123 & new_G3728_;
  assign new_G842_ = new_G3795_ & new_G3815_;
  assign new_G858_ = new_G2500_ & G61 & new_G2476_;
  assign new_G881_ = new_G3737_ & new_G3757_;
  assign new_G4123_ = ~new_G4119_;
  assign new_G4131_ = ~new_G4127_;
  assign new_G4139_ = ~new_G4135_;
  assign new_G4147_ = ~new_G4143_;
  assign new_G4155_ = ~new_G4151_;
  assign new_G4163_ = ~new_G4159_;
  assign new_G4171_ = ~new_G4167_;
  assign new_G4179_ = ~new_G4175_;
  assign new_G4187_ = ~new_G4183_;
  assign new_G4194_ = ~new_G4188_;
  assign new_G4282_ = ~new_G4276_;
  assign new_G4290_ = ~new_G4284_;
  assign new_G4298_ = ~new_G4292_;
  assign new_G4306_ = ~new_G4300_;
  assign new_G4314_ = ~new_G4308_;
  assign new_G4322_ = ~new_G4316_;
  assign new_G4330_ = ~new_G4324_;
  assign new_G4338_ = ~new_G4332_;
  assign new_G4346_ = ~new_G4340_;
  assign new_G1526_ = new_G1697_;
  assign new_G1540_ = ~new_G1528_;
  assign new_G1564_ = ~new_G1552_;
  assign new_G1606_ = new_G1697_;
  assign new_G1621_ = ~new_G1609_;
  assign new_G1645_ = ~new_G1633_;
  assign new_G1661_ = new_G1633_ & G179 & new_G1609_;
  assign new_G1688_ = new_G2826_;
  assign new_G4635_ = ~new_G4631_;
  assign new_G4643_ = ~new_G4639_;
  assign new_G4651_ = ~new_G4647_;
  assign new_G4659_ = ~new_G4655_;
  assign new_G4667_ = ~new_G4663_;
  assign new_G4675_ = ~new_G4671_;
  assign new_G4682_ = ~new_G4676_;
  assign new_G4770_ = ~new_G4764_;
  assign new_G4778_ = ~new_G4772_;
  assign new_G4786_ = ~new_G4780_;
  assign new_G4794_ = ~new_G4788_;
  assign new_G4802_ = ~new_G4796_;
  assign new_G4810_ = ~new_G4804_;
  assign new_G2202_ = new_G1698_;
  assign new_G2215_ = ~new_G2203_;
  assign new_G2238_ = ~new_G2226_;
  assign new_G2279_ = new_G1698_;
  assign new_G2293_ = ~new_G2281_;
  assign new_G2316_ = ~new_G2304_;
  assign new_G2332_ = new_G2304_ & G179 & new_G2281_;
  assign new_G2430_ = ~new_G2418_;
  assign new_G2454_ = ~new_G2442_;
  assign new_G2488_ = ~new_G2476_;
  assign new_G2512_ = ~new_G2500_;
  assign new_G2536_ = ~new_G2533_;
  assign new_G2540_ = ~new_G2537_;
  assign new_G2544_ = ~new_G2541_;
  assign new_G2548_ = ~new_G2545_;
  assign new_G2552_ = ~new_G2549_;
  assign new_G2556_ = ~new_G2553_;
  assign new_G2560_ = ~new_G2557_;
  assign new_G2564_ = ~new_G2561_;
  assign new_G2566_ = new_G2537_ & new_G3553_ & G457;
  assign new_G2572_ = new_G2545_ & new_G3553_ & G468;
  assign new_G2578_ = new_G2553_ & new_G3553_ & G422;
  assign new_G2584_ = new_G2561_ & new_G3553_ & G435;
  assign new_G2590_ = new_G3547_ & new_G2533_;
  assign new_G2595_ = new_G3547_ & new_G2541_;
  assign new_G2600_ = new_G3547_ & new_G2549_;
  assign new_G2605_ = new_G3547_ & new_G2557_;
  assign new_G2630_ = ~new_G2627_;
  assign new_G2634_ = ~new_G2631_;
  assign new_G2638_ = ~new_G2635_;
  assign new_G2642_ = ~new_G2639_;
  assign new_G2646_ = ~new_G2643_;
  assign new_G2650_ = ~new_G2647_;
  assign new_G2654_ = ~new_G2651_;
  assign new_G2658_ = ~new_G2655_;
  assign new_G2660_ = new_G2631_ & new_G3553_ & G389;
  assign new_G2666_ = new_G2639_ & new_G3553_ & G400;
  assign new_G2672_ = new_G2647_ & new_G3553_ & G411;
  assign new_G2678_ = new_G2655_ & new_G3553_ & G374;
  assign new_G2684_ = new_G3547_ & new_G2627_;
  assign new_G2689_ = new_G3547_ & new_G2635_;
  assign new_G2694_ = new_G3547_ & new_G2643_;
  assign new_G2699_ = new_G3547_ & new_G2651_;
  assign new_G2728_ = ~new_G2721_;
  assign new_G2741_ = ~new_G2734_;
  assign new_G2748_ = G292 & new_G2721_;
  assign new_G2750_ = G288 & new_G2721_;
  assign new_G2752_ = G280 & new_G2721_;
  assign new_G2754_ = G272 & new_G2721_;
  assign new_G2756_ = G264 & new_G2721_;
  assign new_G2758_ = G241 & new_G2734_;
  assign new_G2760_ = G233 & new_G2734_;
  assign new_G2762_ = G225 & new_G2734_;
  assign new_G2764_ = G217 & new_G2734_;
  assign new_G2766_ = G209 & new_G2734_;
  assign new_G2827_ = new_G1701_;
  assign new_G2838_ = ~new_G2828_;
  assign new_G2847_ = ~new_G2822_;
  assign new_G2885_ = ~new_G2882_;
  assign new_G2889_ = ~new_G2886_;
  assign new_G2893_ = ~new_G2890_;
  assign new_G2897_ = ~new_G2894_;
  assign new_G2901_ = ~new_G2898_;
  assign new_G2905_ = ~new_G2902_;
  assign new_G2906_ = new_G2393_ & new_G2886_;
  assign new_G2909_ = new_G2894_ & new_G2393_ & G479;
  assign new_G2913_ = new_G2902_ & new_G2393_ & G490;
  assign new_G2918_ = new_G3554_ & new_G2882_;
  assign new_G2922_ = new_G3554_ & new_G2890_;
  assign new_G2927_ = new_G3554_ & new_G2898_;
  assign new_G2951_ = ~new_G2948_;
  assign new_G2955_ = ~new_G2952_;
  assign new_G2959_ = ~new_G2956_;
  assign new_G2963_ = ~new_G2960_;
  assign new_G2967_ = ~new_G2964_;
  assign new_G2971_ = ~new_G2968_;
  assign new_G2973_ = new_G2952_ & new_G3553_ & G503;
  assign new_G2980_ = ~new_G2979_;
  assign new_G2982_ = new_G2960_ & new_G3553_ & G523;
  assign new_G2988_ = new_G2968_ & new_G3553_ & G534;
  assign new_G2994_ = new_G3547_ & new_G2948_;
  assign new_G3001_ = new_G3547_ & new_G2956_;
  assign new_G3006_ = new_G3547_ & new_G2964_;
  assign new_G3027_ = ~new_G3024_;
  assign new_G3031_ = ~new_G3028_;
  assign new_G3035_ = ~new_G3032_;
  assign new_G3039_ = ~new_G3036_;
  assign new_G3043_ = ~new_G3040_;
  assign new_G3047_ = ~new_G3044_;
  assign new_G3051_ = ~new_G3048_;
  assign new_G3055_ = ~new_G3052_;
  assign new_G3056_ = new_G3028_ & new_G2393_ & G389;
  assign new_G3060_ = new_G3036_ & new_G2393_ & G400;
  assign new_G3064_ = new_G3044_ & new_G2393_ & G411;
  assign new_G3068_ = new_G3052_ & new_G2393_ & G374;
  assign new_G3073_ = new_G3554_ & new_G3024_;
  assign new_G3078_ = new_G3554_ & new_G3032_;
  assign new_G3083_ = new_G3554_ & new_G3040_;
  assign new_G3088_ = new_G3554_ & new_G3048_;
  assign new_G3099_ = ~new_G3092_;
  assign new_G3112_ = ~new_G3105_;
  assign new_G3119_ = G372 & new_G3092_;
  assign new_G3121_ = G366 & new_G3092_;
  assign new_G3123_ = G358 & new_G3092_;
  assign new_G3125_ = G348 & new_G3092_;
  assign new_G3126_ = G338 & new_G3092_;
  assign new_G3128_ = G331 & new_G3105_;
  assign new_G3130_ = G323 & new_G3105_;
  assign new_G3132_ = G315 & new_G3105_;
  assign new_G3134_ = G307 & new_G3105_;
  assign new_G3136_ = G299 & new_G3105_;
  assign new_G3187_ = ~new_G3181_;
  assign new_G3193_ = G83 & new_G3181_;
  assign new_G3196_ = G86 & new_G3181_;
  assign new_G3199_ = G88 & new_G3181_;
  assign new_G3202_ = G88 & new_G3181_;
  assign new_G3207_ = ~new_G3204_;
  assign new_G3211_ = ~new_G3208_;
  assign new_G3215_ = ~new_G3212_;
  assign new_G3219_ = ~new_G3216_;
  assign new_G3223_ = ~new_G3220_;
  assign new_G3227_ = ~new_G3224_;
  assign new_G3228_ = new_G3208_ & new_G2405_ & G503;
  assign new_G3232_ = new_G2405_ & G514;
  assign new_G3234_ = new_G3216_ & new_G2405_ & G523;
  assign new_G3238_ = new_G3224_ & new_G2405_ & G534;
  assign new_G3243_ = new_G3555_ & new_G3204_;
  assign new_G3247_ = new_G3555_ | G514;
  assign new_G3249_ = new_G3555_ & new_G3212_;
  assign new_G3253_ = new_G3555_ & new_G3220_;
  assign new_G3259_ = ~new_G3256_;
  assign new_G3263_ = ~new_G3260_;
  assign new_G3267_ = ~new_G3264_;
  assign new_G3271_ = ~new_G3268_;
  assign new_G3275_ = ~new_G3272_;
  assign new_G3279_ = ~new_G3276_;
  assign new_G3280_ = new_G2405_ & new_G3260_;
  assign new_G3283_ = new_G3268_ & new_G2405_ & G479;
  assign new_G3287_ = new_G3276_ & new_G2405_ & G490;
  assign new_G3292_ = new_G3555_ & new_G3256_;
  assign new_G3295_ = new_G3555_ & new_G3264_;
  assign new_G3299_ = new_G3555_ & new_G3272_;
  assign new_G3305_ = ~new_G3302_;
  assign new_G3306_ = new_G2816_;
  assign new_G3310_ = new_G2816_;
  assign new_G3317_ = ~new_G3314_;
  assign new_G3318_ = new_G2816_;
  assign new_G3322_ = new_G2816_;
  assign new_G3326_ = new_G2405_ & new_G3302_;
  assign new_G3333_ = new_G2405_ & new_G3314_;
  assign new_G3357_ = ~new_G3354_;
  assign new_G3361_ = ~new_G3358_;
  assign new_G3365_ = ~new_G3362_;
  assign new_G3369_ = ~new_G3366_;
  assign new_G3373_ = ~new_G3370_;
  assign new_G3377_ = ~new_G3374_;
  assign new_G3381_ = ~new_G3378_;
  assign new_G3385_ = ~new_G3382_;
  assign new_G3386_ = new_G3358_ & new_G2393_ & G457;
  assign new_G3390_ = new_G3366_ & new_G2393_ & G468;
  assign new_G3394_ = new_G3374_ & new_G2393_ & G422;
  assign new_G3398_ = new_G3382_ & new_G2393_ & G435;
  assign new_G3403_ = new_G3554_ & new_G3354_;
  assign new_G3408_ = new_G3554_ & new_G3362_;
  assign new_G3413_ = new_G3554_ & new_G3370_;
  assign new_G3418_ = new_G3554_ & new_G3378_;
  assign new_G5088_ = ~new_G5082_;
  assign new_G5089_ = ~new_G5085_;
  assign new_G5096_ = ~new_G5090_;
  assign new_G5097_ = ~new_G5093_;
  assign new_G3489_ = new_G3440_;
  assign new_G3493_ = new_G3440_;
  assign new_G3570_ = ~new_G3558_;
  assign new_G3594_ = ~new_G3582_;
  assign new_G3622_ = ~new_G3616_;
  assign new_G3632_ = ~new_G3628_;
  assign new_G3637_ = G97 & new_G3616_;
  assign new_G3640_ = G94 & new_G3616_;
  assign new_G3643_ = G97 & new_G3616_;
  assign new_G3646_ = G94 & new_G3616_;
  assign new_G3672_ = ~new_G3660_;
  assign new_G3696_ = ~new_G3684_;
  assign new_G3745_ = ~new_G3737_;
  assign new_G3765_ = ~new_G3757_;
  assign new_G3803_ = ~new_G3795_;
  assign new_G3823_ = ~new_G3815_;
  assign new_G5338_ = ~new_G5332_;
  assign new_G5339_ = ~new_G5335_;
  assign new_G5346_ = ~new_G5340_;
  assign new_G5347_ = ~new_G5343_;
  assign new_G5354_ = ~new_G5348_;
  assign new_G5355_ = ~new_G5351_;
  assign new_G3979_ = ~new_G3972_;
  assign new_G3998_ = ~new_G3991_;
  assign new_G4037_ = ~new_G4030_;
  assign new_G4056_ = ~new_G4049_;
  assign new_G4094_ = new_G4110_;
  assign new_G5104_ = ~new_G5098_;
  assign new_G5105_ = ~new_G5101_;
  assign new_G5114_ = ~new_G5108_;
  assign new_G5115_ = ~new_G5111_;
  assign new_G5362_ = ~new_G5356_;
  assign new_G5363_ = ~new_G5359_;
  assign new_G5366_ = new_G2816_;
  assign new_G5373_ = ~new_G5369_;
  assign G993 = new_G1688_;
  assign G978 = new_G1688_;
  assign G949 = new_G1688_;
  assign G939 = new_G1688_;
  assign new_G2568_ = new_G2540_ & G457 & new_G3551_;
  assign new_G2574_ = new_G2548_ & G468 & new_G3551_;
  assign new_G2580_ = new_G2556_ & G422 & new_G3551_;
  assign new_G2586_ = new_G2564_ & G435 & new_G3551_;
  assign new_G2592_ = new_G3549_ & new_G2536_;
  assign new_G2597_ = new_G3549_ & new_G2544_;
  assign new_G2602_ = new_G3549_ & new_G2552_;
  assign new_G2607_ = new_G3549_ & new_G2560_;
  assign new_G2662_ = new_G2634_ & G389 & new_G3551_;
  assign new_G2668_ = new_G2642_ & G400 & new_G3551_;
  assign new_G2674_ = new_G2650_ & G411 & new_G3551_;
  assign new_G2680_ = new_G2658_ & G374 & new_G3551_;
  assign new_G2686_ = new_G3549_ & new_G2630_;
  assign new_G2691_ = new_G3549_ & new_G2638_;
  assign new_G2696_ = new_G3549_ & new_G2646_;
  assign new_G2701_ = new_G3549_ & new_G2654_;
  assign new_G2907_ = new_G2370_ & new_G2889_;
  assign new_G2910_ = new_G2897_ & G479 & new_G2370_;
  assign new_G2914_ = new_G2905_ & G490 & new_G2370_;
  assign new_G2920_ = new_G3556_ & new_G2885_;
  assign new_G2924_ = new_G3556_ & new_G2893_;
  assign new_G2929_ = new_G3556_ & new_G2901_;
  assign new_G2975_ = new_G2955_ & G503 & new_G3551_;
  assign new_G2984_ = new_G2963_ & G523 & new_G3551_;
  assign new_G2990_ = new_G2971_ & G534 & new_G3551_;
  assign new_G2996_ = new_G3549_ & new_G2951_;
  assign new_G3003_ = new_G3549_ & new_G2959_;
  assign new_G3008_ = new_G3549_ & new_G2967_;
  assign new_G3015_ = new_G2980_ & new_G2999_;
  assign new_G3057_ = new_G3031_ & G389 & new_G2370_;
  assign new_G3061_ = new_G3039_ & G400 & new_G2370_;
  assign new_G3065_ = new_G3047_ & G411 & new_G2370_;
  assign new_G3069_ = new_G3055_ & G374 & new_G2370_;
  assign new_G3075_ = new_G3556_ & new_G3027_;
  assign new_G3080_ = new_G3556_ & new_G3035_;
  assign new_G3085_ = new_G3556_ & new_G3043_;
  assign new_G3090_ = new_G3556_ & new_G3051_;
  assign new_G3229_ = new_G3211_ & G503 & new_G2382_;
  assign new_G3233_ = ~new_G3232_;
  assign new_G3235_ = new_G3219_ & G523 & new_G2382_;
  assign new_G3239_ = new_G3227_ & G534 & new_G2382_;
  assign new_G3244_ = new_G2361_ & new_G3207_;
  assign new_G3250_ = new_G2361_ & new_G3215_;
  assign new_G3254_ = new_G2361_ & new_G3223_;
  assign new_G3281_ = new_G2382_ & new_G3263_;
  assign new_G3284_ = new_G3271_ & G479 & new_G2382_;
  assign new_G3288_ = new_G3279_ & G490 & new_G2382_;
  assign new_G3293_ = new_G2361_ & new_G3259_;
  assign new_G3296_ = new_G2361_ & new_G3267_;
  assign new_G3300_ = new_G2361_ & new_G3275_;
  assign new_G3327_ = new_G2382_ & new_G3305_;
  assign new_G3334_ = new_G2382_ & new_G3317_;
  assign new_G3387_ = new_G3361_ & G457 & new_G2370_;
  assign new_G3391_ = new_G3369_ & G468 & new_G2370_;
  assign new_G3395_ = new_G3377_ & G422 & new_G2370_;
  assign new_G3399_ = new_G3385_ & G435 & new_G2370_;
  assign new_G3405_ = new_G3556_ & new_G3357_;
  assign new_G3410_ = new_G3556_ & new_G3365_;
  assign new_G3415_ = new_G3556_ & new_G3373_;
  assign new_G3420_ = new_G3556_ & new_G3381_;
  assign new_G3422_ = ~new_G5085_ | ~new_G5088_;
  assign new_G3423_ = ~new_G5082_ | ~new_G5089_;
  assign new_G3431_ = ~new_G5093_ | ~new_G5096_;
  assign new_G3432_ = ~new_G5090_ | ~new_G5097_;
  assign new_G3895_ = ~new_G5335_ | ~new_G5338_;
  assign new_G3896_ = ~new_G5332_ | ~new_G5339_;
  assign new_G3904_ = ~new_G5343_ | ~new_G5346_;
  assign new_G3905_ = ~new_G5340_ | ~new_G5347_;
  assign new_G3913_ = ~new_G5351_ | ~new_G5354_;
  assign new_G3914_ = ~new_G5348_ | ~new_G5355_;
  assign G889 = new_G4094_;
  assign new_G5106_ = ~new_G5101_ | ~new_G5104_;
  assign new_G5107_ = ~new_G5098_ | ~new_G5105_;
  assign new_G5116_ = ~new_G5111_ | ~new_G5114_;
  assign new_G5117_ = ~new_G5108_ | ~new_G5115_;
  assign new_G5364_ = ~new_G5359_ | ~new_G5362_;
  assign new_G5365_ = ~new_G5356_ | ~new_G5363_;
  assign G593 = ~new_G4094_;
  assign new_G2880_ = new_G2838_ & new_G2847_;
  assign new_G2881_ = new_G2828_ & new_G2847_;
  assign new_G1579_ = new_G1552_ & G200 & new_G1540_;
  assign new_G1585_ = new_G1552_ & G203 & new_G1540_;
  assign new_G1591_ = new_G1552_ & G197 & new_G1540_;
  assign new_G1597_ = new_G1552_ & G194 & new_G1540_;
  assign new_G1603_ = new_G1552_ & G191 & new_G1540_;
  assign new_G1667_ = new_G1633_ & G182 & new_G1621_;
  assign new_G1673_ = new_G1633_ & G188 & new_G1621_;
  assign new_G1679_ = new_G1633_ & G155 & new_G1621_;
  assign new_G1685_ = new_G1633_ & G149 & new_G1621_;
  assign new_G2876_ = new_G2838_ & new_G2847_;
  assign new_G2877_ = new_G2828_ & new_G2847_;
  assign new_G2253_ = new_G2226_ & G200 & new_G2215_;
  assign new_G2259_ = new_G2226_ & G203 & new_G2215_;
  assign new_G2265_ = new_G2226_ & G197 & new_G2215_;
  assign new_G2271_ = new_G2226_ & G194 & new_G2215_;
  assign new_G2277_ = new_G2226_ & G191 & new_G2215_;
  assign new_G2338_ = new_G2304_ & G182 & new_G2293_;
  assign new_G2344_ = new_G2304_ & G188 & new_G2293_;
  assign new_G2350_ = new_G2304_ & G155 & new_G2293_;
  assign new_G2356_ = new_G2304_ & G149 & new_G2293_;
  assign new_G2868_ = new_G2838_ & new_G2847_;
  assign new_G2869_ = new_G2828_ & new_G2847_;
  assign new_G710_ = new_G3684_ & G109 & new_G3672_;
  assign new_G2872_ = new_G2838_ & new_G2847_;
  assign new_G2873_ = new_G2828_ & new_G2847_;
  assign new_G720_ = new_G2442_ & G11 & new_G2430_;
  assign new_G725_ = new_G3582_ & G109 & new_G3570_;
  assign new_G730_ = new_G3582_ & G46 & new_G3570_;
  assign new_G735_ = new_G3582_ & G100 & new_G3570_;
  assign new_G740_ = new_G3582_ & G91 & new_G3570_;
  assign new_G745_ = new_G3582_ & G43 & new_G3570_;
  assign new_G750_ = new_G2442_ & G76 & new_G2430_;
  assign new_G755_ = new_G2442_ & G73 & new_G2430_;
  assign new_G760_ = new_G2442_ & G67 & new_G2430_;
  assign new_G765_ = new_G2442_ & G14 & new_G2430_;
  assign new_G770_ = new_G3684_ & G46 & new_G3672_;
  assign new_G775_ = new_G3684_ & G100 & new_G3672_;
  assign new_G780_ = new_G3684_ & G91 & new_G3672_;
  assign new_G785_ = new_G3684_ & G43 & new_G3672_;
  assign new_G790_ = new_G2500_ & G76 & new_G2488_;
  assign new_G795_ = new_G2500_ & G73 & new_G2488_;
  assign new_G800_ = new_G2500_ & G67 & new_G2488_;
  assign new_G805_ = new_G2500_ & G14 & new_G2488_;
  assign new_G841_ = new_G3815_ & G120 & new_G3803_;
  assign new_G857_ = new_G2500_ & G11 & new_G2488_;
  assign new_G880_ = new_G3757_ & G118 & new_G3745_;
  assign new_G1660_ = new_G1633_ & G176 & new_G1621_;
  assign new_G2331_ = new_G2304_ & G176 & new_G2293_;
  assign new_G2569_ = new_G2566_ | new_G2568_;
  assign new_G2575_ = new_G2572_ | new_G2574_;
  assign new_G2581_ = new_G2578_ | new_G2580_;
  assign new_G2587_ = new_G2584_ | new_G2586_;
  assign new_G2593_ = G457 | new_G2590_ | new_G2592_;
  assign new_G2598_ = G468 | new_G2595_ | new_G2597_;
  assign new_G2603_ = G422 | new_G2600_ | new_G2602_;
  assign new_G2608_ = G435 | new_G2605_ | new_G2607_;
  assign new_G2663_ = new_G2660_ | new_G2662_;
  assign new_G2669_ = new_G2666_ | new_G2668_;
  assign new_G2675_ = new_G2672_ | new_G2674_;
  assign new_G2681_ = new_G2678_ | new_G2680_;
  assign new_G2687_ = G389 | new_G2684_ | new_G2686_;
  assign new_G2692_ = G400 | new_G2689_ | new_G2691_;
  assign new_G2697_ = G411 | new_G2694_ | new_G2696_;
  assign new_G2702_ = G374 | new_G2699_ | new_G2701_;
  assign new_G2747_ = G289 & new_G2728_;
  assign new_G2749_ = G281 & new_G2728_;
  assign new_G2751_ = G273 & new_G2728_;
  assign new_G2753_ = G265 & new_G2728_;
  assign new_G2755_ = G257 & new_G2728_;
  assign new_G2757_ = G234 & new_G2741_;
  assign new_G2759_ = G226 & new_G2741_;
  assign new_G2761_ = G218 & new_G2741_;
  assign new_G2763_ = G210 & new_G2741_;
  assign new_G2765_ = G206 & new_G2741_;
  assign new_G2857_ = ~new_G2847_;
  assign new_G2908_ = new_G2906_ | new_G2907_;
  assign new_G2911_ = new_G2909_ | new_G2910_;
  assign new_G2915_ = new_G2913_ | new_G2914_;
  assign new_G2925_ = G479 | new_G2922_ | new_G2924_;
  assign new_G2930_ = G490 | new_G2927_ | new_G2929_;
  assign new_G2933_ = new_G2918_ | new_G2920_;
  assign new_G2976_ = new_G2973_ | new_G2975_;
  assign new_G2985_ = new_G2982_ | new_G2984_;
  assign new_G2991_ = new_G2988_ | new_G2990_;
  assign new_G2997_ = G503 | new_G2994_ | new_G2996_;
  assign new_G3004_ = G523 | new_G3001_ | new_G3003_;
  assign new_G3009_ = G534 | new_G3006_ | new_G3008_;
  assign new_G3058_ = new_G3056_ | new_G3057_;
  assign new_G3062_ = new_G3060_ | new_G3061_;
  assign new_G3066_ = new_G3064_ | new_G3065_;
  assign new_G3070_ = new_G3068_ | new_G3069_;
  assign new_G3076_ = G389 | new_G3073_ | new_G3075_;
  assign new_G3081_ = G400 | new_G3078_ | new_G3080_;
  assign new_G3086_ = G411 | new_G3083_ | new_G3085_;
  assign new_G3091_ = G374 | new_G3088_ | new_G3090_;
  assign new_G3118_ = G369 & new_G3099_;
  assign new_G3120_ = G361 & new_G3099_;
  assign new_G3122_ = G351 & new_G3099_;
  assign new_G3124_ = G341 & new_G3099_;
  assign new_G3127_ = G324 & new_G3112_;
  assign new_G3129_ = G316 & new_G3112_;
  assign new_G3131_ = G308 & new_G3112_;
  assign new_G3133_ = G302 & new_G3112_;
  assign new_G3135_ = G293 & new_G3112_;
  assign new_G3147_ = new_G3099_ | new_G3126_;
  assign new_G3192_ = G83 & new_G3187_;
  assign new_G3195_ = G87 & new_G3187_;
  assign new_G3198_ = G34 & new_G3187_;
  assign new_G3201_ = G34 & new_G3187_;
  assign new_G3230_ = new_G3228_ | new_G3229_;
  assign new_G3236_ = new_G3234_ | new_G3235_;
  assign new_G3240_ = new_G3238_ | new_G3239_;
  assign new_G3245_ = G503 | new_G3243_ | new_G3244_;
  assign new_G3251_ = G523 | new_G3249_ | new_G3250_;
  assign new_G3255_ = G534 | new_G3253_ | new_G3254_;
  assign new_G3282_ = new_G3280_ | new_G3281_;
  assign new_G3285_ = new_G3283_ | new_G3284_;
  assign new_G3289_ = new_G3287_ | new_G3288_;
  assign new_G3297_ = G479 | new_G3295_ | new_G3296_;
  assign new_G3301_ = G490 | new_G3299_ | new_G3300_;
  assign new_G3309_ = ~new_G3306_;
  assign new_G3313_ = ~new_G3310_;
  assign new_G3321_ = ~new_G3318_;
  assign new_G3325_ = ~new_G3322_;
  assign new_G3328_ = new_G3326_ | new_G3327_;
  assign new_G3329_ = new_G3310_ & new_G2405_ & G446;
  assign new_G3335_ = new_G3333_ | new_G3334_;
  assign new_G3336_ = new_G3322_ & new_G2405_ & G446;
  assign new_G3341_ = new_G3555_ & new_G3306_;
  assign new_G3345_ = new_G3555_ & new_G3318_;
  assign new_G3388_ = new_G3386_ | new_G3387_;
  assign new_G3392_ = new_G3390_ | new_G3391_;
  assign new_G3396_ = new_G3394_ | new_G3395_;
  assign new_G3400_ = new_G3398_ | new_G3399_;
  assign new_G3406_ = G457 | new_G3403_ | new_G3405_;
  assign new_G3411_ = G468 | new_G3408_ | new_G3410_;
  assign new_G3416_ = G422 | new_G3413_ | new_G3415_;
  assign new_G3421_ = G435 | new_G3418_ | new_G3420_;
  assign new_G3424_ = ~new_G3422_ | ~new_G3423_;
  assign new_G3433_ = ~new_G3431_ | ~new_G3432_;
  assign new_G3492_ = ~new_G3489_;
  assign new_G3496_ = ~new_G3493_;
  assign new_G3780_ = new_G3757_ & G117 & new_G3745_;
  assign new_G3783_ = new_G3757_ & G126 & new_G3745_;
  assign new_G3786_ = new_G3757_ & G127 & new_G3745_;
  assign new_G3789_ = new_G3757_ & G128 & new_G3745_;
  assign new_G3838_ = new_G3815_ & G131 & new_G3803_;
  assign new_G3841_ = new_G3815_ & G129 & new_G3803_;
  assign new_G3844_ = new_G3815_ & G119 & new_G3803_;
  assign new_G3847_ = new_G3815_ & G130 & new_G3803_;
  assign new_G3897_ = ~new_G3895_ | ~new_G3896_;
  assign new_G3906_ = ~new_G3904_ | ~new_G3905_;
  assign new_G3915_ = ~new_G3913_ | ~new_G3914_;
  assign new_G4011_ = new_G3991_ & G122 & new_G3979_;
  assign new_G4014_ = new_G3991_ & G113 & new_G3979_;
  assign new_G4017_ = new_G3991_ & G53 & new_G3979_;
  assign new_G4020_ = new_G3991_ & G114 & new_G3979_;
  assign new_G4023_ = new_G3991_ & G115 & new_G3979_;
  assign new_G4069_ = new_G4049_ & G52 & new_G4037_;
  assign new_G4072_ = new_G4049_ & G112 & new_G4037_;
  assign new_G4075_ = new_G4049_ & G116 & new_G4037_;
  assign new_G4078_ = new_G4049_ & G121 & new_G4037_;
  assign new_G4081_ = new_G4049_ & G123 & new_G4037_;
  assign new_G5206_ = ~new_G5116_ | ~new_G5117_;
  assign new_G5209_ = ~new_G5106_ | ~new_G5107_;
  assign new_G5307_ = new_G3233_ & new_G3247_;
  assign new_G5322_ = new_G3292_ | new_G3293_;
  assign new_G5372_ = ~new_G5366_;
  assign new_G5375_ = ~new_G5366_ | ~new_G5373_;
  assign new_G5399_ = ~new_G5364_ | ~new_G5365_;
  assign new_G2813_ = ~new_G3015_;
  assign new_G3197_ = new_G3195_ | new_G3196_;
  assign new_G3200_ = new_G3198_ | new_G3199_;
  assign new_G3203_ = new_G3201_ | new_G3202_;
  assign new_G3194_ = new_G3192_ | new_G3193_;
  assign new_G2570_ = ~new_G2569_;
  assign new_G2576_ = ~new_G2575_;
  assign new_G2582_ = ~new_G2581_;
  assign new_G2588_ = ~new_G2587_;
  assign new_G2664_ = ~new_G2663_;
  assign new_G2670_ = ~new_G2669_;
  assign new_G2676_ = ~new_G2675_;
  assign new_G2682_ = ~new_G2681_;
  assign new_G2767_ = new_G2749_ | new_G2750_;
  assign new_G2772_ = new_G2751_ | new_G2752_;
  assign new_G2776_ = new_G2753_ | new_G2754_;
  assign new_G2780_ = new_G2755_ | new_G2756_;
  assign new_G2784_ = new_G2757_ | new_G2758_;
  assign new_G2788_ = new_G2759_ | new_G2760_;
  assign new_G2794_ = new_G2761_ | new_G2762_;
  assign new_G2798_ = new_G2763_ | new_G2764_;
  assign new_G2802_ = new_G2765_ | new_G2766_;
  assign new_G2912_ = ~new_G2911_;
  assign new_G2916_ = ~new_G2915_;
  assign new_G2936_ = ~new_G2908_;
  assign new_G2977_ = ~new_G2976_;
  assign new_G2986_ = ~new_G2985_;
  assign new_G2992_ = ~new_G2991_;
  assign new_G3059_ = ~new_G3058_;
  assign new_G3063_ = ~new_G3062_;
  assign new_G3067_ = ~new_G3066_;
  assign new_G3071_ = ~new_G3070_;
  assign new_G3137_ = new_G3120_ | new_G3121_;
  assign new_G3139_ = new_G3122_ | new_G3123_;
  assign new_G3143_ = new_G3124_ | new_G3125_;
  assign new_G3151_ = new_G3127_ | new_G3128_;
  assign new_G3155_ = new_G3129_ | new_G3130_;
  assign new_G3161_ = new_G3131_ | new_G3132_;
  assign new_G3165_ = new_G3133_ | new_G3134_;
  assign new_G3167_ = new_G3135_ | new_G3136_;
  assign new_G3231_ = ~new_G3230_;
  assign new_G3237_ = ~new_G3236_;
  assign new_G3241_ = ~new_G3240_;
  assign new_G3286_ = ~new_G3285_;
  assign new_G3290_ = ~new_G3289_;
  assign new_G3330_ = new_G3313_ & G446 & new_G2382_;
  assign new_G3337_ = new_G3325_ & G446 & new_G2382_;
  assign new_G3342_ = new_G2361_ & new_G3309_;
  assign new_G3346_ = new_G2361_ & new_G3321_;
  assign new_G3348_ = ~new_G3328_;
  assign new_G3352_ = ~new_G3335_;
  assign new_G3389_ = ~new_G3388_;
  assign new_G3393_ = ~new_G3392_;
  assign new_G3397_ = ~new_G3396_;
  assign new_G3401_ = ~new_G3400_;
  assign new_G3845_ = new_G3823_ & new_G3015_ & new_G3803_;
  assign new_G5126_ = new_G3118_ | new_G3119_;
  assign new_G5178_ = new_G2747_ | new_G2748_;
  assign new_G5325_ = ~new_G3282_;
  assign new_G5374_ = ~new_G5369_ | ~new_G5372_;
  assign new_G2810_ = ~new_G2933_;
  assign new_G635_ = new_G3197_ & new_G3176_;
  assign new_G2878_ = new_G2857_ & G24 & new_G2838_;
  assign new_G2879_ = new_G2857_ & G25 & new_G2828_;
  assign new_G2874_ = new_G2857_ & G26 & new_G2838_;
  assign new_G2875_ = new_G2857_ & G81 & new_G2828_;
  assign new_G703_ = new_G3200_ & new_G3176_;
  assign new_G2866_ = new_G2857_ & G79 & new_G2838_;
  assign new_G2867_ = new_G2857_ & G23 & new_G2828_;
  assign new_G2870_ = new_G2857_ & G82 & new_G2838_;
  assign new_G2871_ = new_G2857_ & G80 & new_G2828_;
  assign new_G716_ = new_G3203_ & new_G3176_;
  assign new_G819_ = new_G3194_ & new_G3176_;
  assign new_G1789_ = new_G3147_ & G514;
  assign new_G2036_ = G514 & new_G3147_;
  assign new_G2611_ = new_G2570_ & new_G2593_;
  assign new_G2615_ = new_G2576_ & new_G2598_;
  assign new_G2619_ = new_G2582_ & new_G2603_;
  assign new_G2623_ = new_G2588_ & new_G2608_;
  assign new_G2705_ = new_G2664_ & new_G2687_;
  assign new_G2709_ = new_G2670_ & new_G2692_;
  assign new_G2713_ = new_G2676_ & new_G2697_;
  assign new_G2717_ = new_G2682_ & new_G2702_;
  assign new_G2939_ = new_G2912_ & new_G2925_;
  assign new_G2942_ = new_G2916_ & new_G2930_;
  assign new_G2945_ = new_G2933_;
  assign new_G3012_ = new_G2977_ & new_G2997_;
  assign new_G3018_ = new_G2986_ & new_G3004_;
  assign new_G3021_ = new_G2992_ & new_G3009_;
  assign new_G3331_ = new_G3329_ | new_G3330_;
  assign new_G3338_ = new_G3336_ | new_G3337_;
  assign new_G3343_ = G446 | new_G3341_ | new_G3342_;
  assign new_G3347_ = G446 | new_G3345_ | new_G3346_;
  assign new_G3428_ = ~new_G3424_;
  assign new_G3437_ = ~new_G3433_;
  assign new_G3514_ = new_G3489_ & new_G3433_ & new_G3424_;
  assign new_G3836_ = new_G3823_ & new_G3352_ & new_G3803_;
  assign new_G3852_ = new_G3071_ & new_G3091_;
  assign new_G5311_ = ~new_G5307_;
  assign new_G3901_ = ~new_G3897_;
  assign new_G3910_ = ~new_G3906_;
  assign new_G3934_ = new_G3915_;
  assign new_G3938_ = new_G3915_;
  assign new_G4652_ = new_G3147_;
  assign new_G4783_ = new_G3147_;
  assign new_G5137_ = new_G3147_;
  assign new_G5212_ = ~new_G5206_;
  assign new_G5213_ = ~new_G5209_;
  assign new_G5260_ = new_G3063_ & new_G3081_;
  assign new_G5263_ = new_G3067_ & new_G3086_;
  assign new_G5268_ = new_G3401_ & new_G3421_;
  assign new_G5271_ = new_G3059_ & new_G3076_;
  assign new_G5276_ = new_G3393_ & new_G3411_;
  assign new_G5279_ = new_G3397_ & new_G3416_;
  assign new_G5289_ = new_G3389_ & new_G3406_;
  assign new_G5296_ = new_G3237_ & new_G3251_;
  assign new_G5299_ = new_G3241_ & new_G3255_;
  assign new_G5304_ = new_G3231_ & new_G3245_;
  assign new_G5312_ = new_G3286_ & new_G3297_;
  assign new_G5315_ = new_G3290_ & new_G3301_;
  assign new_G5328_ = ~new_G5322_;
  assign new_G5396_ = ~new_G5374_ | ~new_G5375_;
  assign new_G5403_ = ~new_G5399_;
  assign new_G1286_ = G446 & new_G2802_;
  assign new_G2809_ = ~new_G2936_;
  assign new_G597_ = ~new_G3348_;
  assign new_G1031_ = new_G2802_ & G446;
  assign G636 = ~new_G635_;
  assign new_G637_ = new_G2881_ | new_G2880_ | new_G2878_ | new_G2879_;
  assign new_G671_ = new_G2877_ | new_G2876_ | new_G2874_ | new_G2875_;
  assign G704 = ~new_G703_;
  assign new_G705_ = new_G2869_ | new_G2868_ | new_G2866_ | new_G2867_;
  assign new_G713_ = new_G2873_ | new_G2872_ | new_G2870_ | new_G2871_;
  assign G717 = ~new_G716_;
  assign G820 = ~new_G819_;
  assign new_G1046_ = new_G2798_ & G457;
  assign new_G1064_ = new_G2794_ & G468;
  assign new_G1071_ = G422 & new_G2788_;
  assign new_G1097_ = new_G2784_ & G435;
  assign new_G1111_ = new_G2780_ & G389;
  assign new_G1128_ = new_G2776_ & G400;
  assign new_G1145_ = new_G2772_ & G411;
  assign new_G1160_ = new_G2767_ & G374;
  assign new_G1301_ = G457 & new_G2798_;
  assign new_G1318_ = G468 & new_G2794_;
  assign new_G1324_ = G422 & new_G2788_;
  assign new_G1341_ = G435 & new_G2784_;
  assign new_G1359_ = G389 & new_G2780_;
  assign new_G1382_ = G400 & new_G2776_;
  assign new_G1404_ = G411 & new_G2772_;
  assign new_G1412_ = G374 & new_G2767_;
  assign new_G1704_ = ~new_G3167_;
  assign new_G1712_ = ~new_G3165_;
  assign new_G1724_ = new_G3165_;
  assign new_G1742_ = new_G3161_ & G479;
  assign new_G1749_ = G490 & new_G3155_;
  assign new_G1775_ = new_G3151_ & G503;
  assign new_G1806_ = new_G3143_ & G523;
  assign new_G1823_ = new_G3139_ & G534;
  assign new_G1829_ = ~new_G3137_;
  assign new_G1837_ = new_G3137_;
  assign new_G1958_ = ~new_G3167_;
  assign new_G1966_ = ~new_G3165_;
  assign new_G1978_ = new_G3165_;
  assign new_G1995_ = G479 & new_G3161_;
  assign new_G2001_ = G490 & new_G3155_;
  assign new_G2018_ = G503 & new_G3151_;
  assign new_G2059_ = G523 & new_G3143_;
  assign new_G2081_ = G534 & new_G3139_;
  assign new_G2089_ = new_G3137_;
  assign new_G2106_ = ~new_G3137_;
  assign new_G3170_ = new_G3167_;
  assign new_G3332_ = ~new_G3331_;
  assign new_G3339_ = ~new_G3338_;
  assign new_G5132_ = ~new_G5126_;
  assign new_G5184_ = ~new_G5178_;
  assign new_G3853_ = ~new_G3852_;
  assign new_G3874_ = ~new_G3348_;
  assign new_G4076_ = new_G4056_ & new_G2936_ & new_G4037_;
  assign new_G4116_ = new_G2802_;
  assign new_G4124_ = new_G2798_;
  assign new_G4132_ = new_G2794_;
  assign new_G4140_ = new_G2788_;
  assign new_G4148_ = new_G2784_;
  assign new_G4156_ = new_G2780_;
  assign new_G4164_ = new_G2776_;
  assign new_G4172_ = new_G2772_;
  assign new_G4180_ = new_G2767_;
  assign new_G4228_ = ~G422 & ~new_G2788_;
  assign new_G4279_ = new_G2802_;
  assign new_G4287_ = new_G2798_;
  assign new_G4295_ = new_G2794_;
  assign new_G4303_ = new_G2784_;
  assign new_G4311_ = new_G2780_;
  assign new_G4319_ = new_G2776_;
  assign new_G4327_ = new_G2772_;
  assign new_G4335_ = new_G2788_;
  assign new_G4343_ = new_G2767_;
  assign new_G4348_ = ~G422 & ~new_G2788_;
  assign new_G4464_ = ~G374 & ~new_G2767_;
  assign new_G4628_ = new_G3161_;
  assign new_G4636_ = new_G3155_;
  assign new_G4644_ = new_G3151_;
  assign new_G4660_ = new_G3143_;
  assign new_G4668_ = new_G3139_;
  assign new_G4716_ = ~G490 & ~new_G3155_;
  assign new_G4767_ = new_G3161_;
  assign new_G4775_ = new_G3151_;
  assign new_G4791_ = new_G3143_;
  assign new_G4799_ = new_G3139_;
  assign new_G4807_ = new_G3155_;
  assign new_G4812_ = ~G490 & ~new_G3155_;
  assign new_G5118_ = new_G3139_;
  assign new_G5121_ = new_G3143_;
  assign new_G5129_ = new_G3137_;
  assign new_G5134_ = new_G3151_;
  assign new_G5142_ = new_G3161_;
  assign new_G5145_ = new_G3155_;
  assign new_G5152_ = new_G3167_;
  assign new_G5155_ = new_G3165_;
  assign new_G5162_ = new_G2788_;
  assign new_G5165_ = new_G2784_;
  assign new_G5170_ = new_G2798_;
  assign new_G5173_ = new_G2794_;
  assign new_G5181_ = new_G2802_;
  assign new_G5186_ = new_G2772_;
  assign new_G5189_ = new_G2767_;
  assign new_G5196_ = new_G2780_;
  assign new_G5199_ = new_G2776_;
  assign new_G5214_ = ~new_G5209_ | ~new_G5212_;
  assign new_G5215_ = ~new_G5206_ | ~new_G5213_;
  assign new_G5329_ = ~new_G5325_;
  assign new_G5330_ = ~new_G5325_ | ~new_G5328_;
  assign new_G2807_ = ~new_G2942_;
  assign new_G2808_ = ~new_G2939_;
  assign new_G2811_ = ~new_G3021_;
  assign new_G2812_ = ~new_G3018_;
  assign new_G2814_ = ~new_G3012_;
  assign new_G2626_ = ~new_G2623_;
  assign new_G2622_ = ~new_G2619_;
  assign new_G2618_ = ~new_G2615_;
  assign new_G2614_ = ~new_G2611_;
  assign new_G2720_ = ~new_G2717_;
  assign new_G2716_ = ~new_G2713_;
  assign new_G2712_ = ~new_G2709_;
  assign new_G2708_ = ~new_G2705_;
  assign G639 = new_G637_ & new_G2827_;
  assign G673 = new_G671_ & new_G2827_;
  assign G707 = new_G705_ & new_G2827_;
  assign G715 = new_G713_ & new_G2827_;
  assign new_G3731_ = new_G3721_ & new_G2945_ & new_G3728_;
  assign new_G4658_ = ~new_G4652_;
  assign new_G1777_ = ~new_G4652_ | ~new_G4659_;
  assign new_G2019_ = ~new_G4783_ | ~new_G4786_;
  assign new_G4787_ = ~new_G4783_;
  assign new_G3350_ = new_G3332_ & new_G3343_;
  assign new_G3353_ = new_G3339_ & new_G3347_;
  assign new_G5141_ = ~new_G5137_;
  assign new_G3513_ = new_G3492_ & new_G3428_ & new_G3433_;
  assign new_G3516_ = new_G3496_ & new_G3424_ & new_G3437_;
  assign new_G3517_ = new_G3493_ & new_G3437_ & new_G3428_;
  assign new_G3778_ = new_G3765_ & new_G2717_ & new_G3745_;
  assign new_G3781_ = new_G3765_ & new_G2713_ & new_G3745_;
  assign new_G3784_ = new_G3765_ & new_G2709_ & new_G3745_;
  assign new_G3787_ = new_G3765_ & new_G2705_ & new_G3745_;
  assign new_G3839_ = new_G3823_ & new_G3021_ & new_G3803_;
  assign new_G3842_ = new_G3823_ & new_G3018_ & new_G3803_;
  assign new_G5266_ = ~new_G5260_;
  assign new_G5267_ = ~new_G5263_;
  assign new_G5274_ = ~new_G5268_;
  assign new_G5275_ = ~new_G5271_;
  assign new_G5302_ = ~new_G5296_;
  assign new_G5303_ = ~new_G5299_;
  assign new_G5310_ = ~new_G5304_;
  assign new_G3891_ = ~new_G5304_ | ~new_G5311_;
  assign new_G3937_ = ~new_G3934_;
  assign new_G3941_ = ~new_G3938_;
  assign new_G3955_ = new_G3934_ & new_G3906_ & new_G3897_;
  assign new_G3958_ = new_G3938_ & new_G3910_ & new_G3901_;
  assign new_G4009_ = new_G3998_ & new_G2623_ & new_G3979_;
  assign new_G4012_ = new_G3998_ & new_G2619_ & new_G3979_;
  assign new_G4015_ = new_G3998_ & new_G2615_ & new_G3979_;
  assign new_G4018_ = new_G3998_ & new_G2611_ & new_G3979_;
  assign new_G4067_ = new_G4056_ & new_G3012_ & new_G4037_;
  assign new_G4070_ = new_G4056_ & new_G2942_ & new_G4037_;
  assign new_G4073_ = new_G4056_ & new_G2939_ & new_G4037_;
  assign new_G4079_ = new_G4056_ & new_G2945_ & new_G4037_;
  assign new_G5239_ = ~new_G5214_ | ~new_G5215_;
  assign new_G5282_ = ~new_G5276_;
  assign new_G5283_ = ~new_G5279_;
  assign new_G5293_ = ~new_G5289_;
  assign new_G5318_ = ~new_G5312_;
  assign new_G5319_ = ~new_G5315_;
  assign new_G5331_ = ~new_G5322_ | ~new_G5329_;
  assign new_G5402_ = ~new_G5396_;
  assign new_G5405_ = ~new_G5396_ | ~new_G5403_;
  assign new_G595_ = new_G2810_ & new_G2809_ & new_G2807_ & new_G2808_;
  assign new_G596_ = new_G2814_ & new_G2813_ & new_G2811_ & new_G2812_;
  assign new_G607_ = new_G2614_ & new_G2618_ & new_G2626_ & new_G2622_;
  assign new_G608_ = new_G2708_ & new_G2712_ & new_G2720_ & new_G2716_;
  assign new_G1845_ = new_G1704_ & new_G1724_;
  assign new_G1846_ = new_G1742_ & new_G1712_ & new_G1704_;
  assign new_G2115_ = new_G1958_ & new_G1978_;
  assign new_G2116_ = new_G1995_ & new_G1966_ & new_G1958_;
  assign new_G4122_ = ~new_G4116_;
  assign new_G1022_ = ~new_G4116_ | ~new_G4123_;
  assign new_G4130_ = ~new_G4124_;
  assign new_G1033_ = ~new_G4124_ | ~new_G4131_;
  assign new_G4138_ = ~new_G4132_;
  assign new_G1051_ = ~new_G4132_ | ~new_G4139_;
  assign new_G4146_ = ~new_G4140_;
  assign new_G1079_ = ~new_G4140_ | ~new_G4147_;
  assign new_G4154_ = ~new_G4148_;
  assign new_G1088_ = ~new_G4148_ | ~new_G4155_;
  assign new_G4162_ = ~new_G4156_;
  assign new_G1099_ = ~new_G4156_ | ~new_G4163_;
  assign new_G4170_ = ~new_G4164_;
  assign new_G1115_ = ~new_G4164_ | ~new_G4171_;
  assign new_G4178_ = ~new_G4172_;
  assign new_G1133_ = ~new_G4172_ | ~new_G4179_;
  assign new_G4186_ = ~new_G4180_;
  assign new_G1151_ = ~new_G4180_ | ~new_G4187_;
  assign new_G4234_ = ~new_G4228_;
  assign new_G1276_ = ~new_G4279_ | ~new_G4282_;
  assign new_G4283_ = ~new_G4279_;
  assign new_G1287_ = ~new_G4287_ | ~new_G4290_;
  assign new_G4291_ = ~new_G4287_;
  assign new_G1305_ = ~new_G4295_ | ~new_G4298_;
  assign new_G4299_ = ~new_G4295_;
  assign new_G1330_ = ~new_G4303_ | ~new_G4306_;
  assign new_G4307_ = ~new_G4303_;
  assign new_G1342_ = ~new_G4311_ | ~new_G4314_;
  assign new_G4315_ = ~new_G4311_;
  assign new_G1363_ = ~new_G4319_ | ~new_G4322_;
  assign new_G4323_ = ~new_G4319_;
  assign new_G1388_ = ~new_G4327_ | ~new_G4330_;
  assign new_G4331_ = ~new_G4327_;
  assign new_G1420_ = ~new_G4335_ | ~new_G4338_;
  assign new_G4339_ = ~new_G4335_;
  assign new_G1428_ = ~new_G4343_ | ~new_G4346_;
  assign new_G4347_ = ~new_G4343_;
  assign new_G4634_ = ~new_G4628_;
  assign new_G1729_ = ~new_G4628_ | ~new_G4635_;
  assign new_G4642_ = ~new_G4636_;
  assign new_G1757_ = ~new_G4636_ | ~new_G4643_;
  assign new_G4650_ = ~new_G4644_;
  assign new_G1766_ = ~new_G4644_ | ~new_G4651_;
  assign new_G1776_ = ~new_G4655_ | ~new_G4658_;
  assign new_G4666_ = ~new_G4660_;
  assign new_G1793_ = ~new_G4660_ | ~new_G4667_;
  assign new_G4674_ = ~new_G4668_;
  assign new_G1811_ = ~new_G4668_ | ~new_G4675_;
  assign new_G1849_ = new_G1712_ & new_G1742_;
  assign new_G1852_ = new_G1712_ & new_G1742_;
  assign new_G1875_ = G54 & new_G1829_;
  assign new_G4722_ = ~new_G4716_;
  assign new_G1982_ = ~new_G4767_ | ~new_G4770_;
  assign new_G4771_ = ~new_G4767_;
  assign new_G2007_ = ~new_G4775_ | ~new_G4778_;
  assign new_G4779_ = ~new_G4775_;
  assign new_G2020_ = ~new_G4780_ | ~new_G4787_;
  assign new_G2040_ = ~new_G4791_ | ~new_G4794_;
  assign new_G4795_ = ~new_G4791_;
  assign new_G2065_ = ~new_G4799_ | ~new_G4802_;
  assign new_G4803_ = ~new_G4799_;
  assign new_G2097_ = ~new_G4807_ | ~new_G4810_;
  assign new_G4811_ = ~new_G4807_;
  assign new_G2119_ = new_G1966_ & new_G1995_;
  assign new_G2122_ = new_G1966_ & new_G1995_;
  assign new_G5124_ = ~new_G5118_;
  assign new_G5125_ = ~new_G5121_;
  assign new_G3452_ = ~new_G5129_ | ~new_G5132_;
  assign new_G5133_ = ~new_G5129_;
  assign new_G5140_ = ~new_G5134_;
  assign new_G3462_ = ~new_G5134_ | ~new_G5141_;
  assign new_G5168_ = ~new_G5162_;
  assign new_G5169_ = ~new_G5165_;
  assign new_G5176_ = ~new_G5170_;
  assign new_G5177_ = ~new_G5173_;
  assign new_G3484_ = ~new_G5181_ | ~new_G5184_;
  assign new_G5185_ = ~new_G5181_;
  assign new_G3515_ = ~new_G3513_ & ~new_G3514_;
  assign new_G3518_ = ~new_G3516_ & ~new_G3517_;
  assign new_G3857_ = ~new_G3853_;
  assign new_G3860_ = ~new_G5263_ | ~new_G5266_;
  assign new_G3861_ = ~new_G5260_ | ~new_G5267_;
  assign new_G3869_ = ~new_G5271_ | ~new_G5274_;
  assign new_G3870_ = ~new_G5268_ | ~new_G5275_;
  assign new_G3878_ = ~new_G3874_;
  assign new_G3881_ = ~new_G5299_ | ~new_G5302_;
  assign new_G3882_ = ~new_G5296_ | ~new_G5303_;
  assign new_G3890_ = ~new_G5307_ | ~new_G5310_;
  assign new_G3954_ = new_G3937_ & new_G3901_ & new_G3906_;
  assign new_G3957_ = new_G3941_ & new_G3897_ & new_G3910_;
  assign new_G4021_ = new_G3998_ & new_G3353_ & new_G3979_;
  assign new_G4099_ = ~new_G3170_;
  assign new_G4236_ = new_G1071_;
  assign new_G4354_ = ~new_G4348_;
  assign new_G4406_ = new_G1324_;
  assign new_G4470_ = ~new_G4464_;
  assign new_G4552_ = new_G1412_;
  assign new_G4679_ = new_G1829_;
  assign new_G4687_ = new_G1704_;
  assign new_G4695_ = new_G1704_;
  assign new_G4703_ = new_G1712_;
  assign new_G4711_ = new_G1712_;
  assign new_G4724_ = new_G1749_;
  assign new_G4818_ = ~new_G4812_;
  assign new_G4855_ = new_G1958_;
  assign new_G4865_ = new_G1966_;
  assign new_G4870_ = new_G2001_;
  assign new_G4913_ = new_G1958_;
  assign new_G4923_ = new_G1966_;
  assign new_G4951_ = new_G2106_;
  assign new_G5006_ = new_G2089_;
  assign new_G5039_ = new_G2106_;
  assign new_G5148_ = ~new_G5142_;
  assign new_G5149_ = ~new_G5145_;
  assign new_G5158_ = ~new_G5152_;
  assign new_G5159_ = ~new_G5155_;
  assign new_G5192_ = ~new_G5186_;
  assign new_G5193_ = ~new_G5189_;
  assign new_G5202_ = ~new_G5196_;
  assign new_G5203_ = ~new_G5199_;
  assign new_G5284_ = ~new_G5279_ | ~new_G5282_;
  assign new_G5285_ = ~new_G5276_ | ~new_G5283_;
  assign new_G5320_ = ~new_G5315_ | ~new_G5318_;
  assign new_G5321_ = ~new_G5312_ | ~new_G5319_;
  assign new_G5386_ = ~new_G5330_ | ~new_G5331_;
  assign new_G5404_ = ~new_G5399_ | ~new_G5402_;
  assign G598 = new_G597_ & new_G595_ & new_G596_;
  assign new_G609_ = ~new_G3350_;
  assign new_G1021_ = ~new_G4119_ | ~new_G4122_;
  assign new_G1032_ = ~new_G4127_ | ~new_G4130_;
  assign new_G1050_ = ~new_G4135_ | ~new_G4138_;
  assign new_G1078_ = ~new_G4143_ | ~new_G4146_;
  assign new_G1087_ = ~new_G4151_ | ~new_G4154_;
  assign new_G1098_ = ~new_G4159_ | ~new_G4162_;
  assign new_G1114_ = ~new_G4167_ | ~new_G4170_;
  assign new_G1132_ = ~new_G4175_ | ~new_G4178_;
  assign new_G1150_ = ~new_G4183_ | ~new_G4186_;
  assign new_G1277_ = ~new_G4276_ | ~new_G4283_;
  assign new_G1288_ = ~new_G4284_ | ~new_G4291_;
  assign new_G1306_ = ~new_G4292_ | ~new_G4299_;
  assign new_G1331_ = ~new_G4300_ | ~new_G4307_;
  assign new_G1343_ = ~new_G4308_ | ~new_G4315_;
  assign new_G1364_ = ~new_G4316_ | ~new_G4323_;
  assign new_G1389_ = ~new_G4324_ | ~new_G4331_;
  assign new_G1421_ = ~new_G4332_ | ~new_G4339_;
  assign new_G1429_ = ~new_G4340_ | ~new_G4347_;
  assign new_G1728_ = ~new_G4631_ | ~new_G4634_;
  assign new_G1756_ = ~new_G4639_ | ~new_G4642_;
  assign new_G1765_ = ~new_G4647_ | ~new_G4650_;
  assign new_G1778_ = ~new_G1776_ | ~new_G1777_;
  assign new_G1792_ = ~new_G4663_ | ~new_G4666_;
  assign new_G1810_ = ~new_G4671_ | ~new_G4674_;
  assign new_G1983_ = ~new_G4764_ | ~new_G4771_;
  assign new_G2008_ = ~new_G4772_ | ~new_G4779_;
  assign new_G2021_ = ~new_G2019_ | ~new_G2020_;
  assign new_G2041_ = ~new_G4788_ | ~new_G4795_;
  assign new_G2066_ = ~new_G4796_ | ~new_G4803_;
  assign new_G2098_ = ~new_G4804_ | ~new_G4811_;
  assign new_G3443_ = ~new_G5121_ | ~new_G5124_;
  assign new_G3444_ = ~new_G5118_ | ~new_G5125_;
  assign new_G3453_ = ~new_G5126_ | ~new_G5133_;
  assign new_G3461_ = ~new_G5137_ | ~new_G5140_;
  assign new_G3466_ = ~new_G5165_ | ~new_G5168_;
  assign new_G3467_ = ~new_G5162_ | ~new_G5169_;
  assign new_G3475_ = ~new_G5173_ | ~new_G5176_;
  assign new_G3476_ = ~new_G5170_ | ~new_G5177_;
  assign new_G3485_ = ~new_G5178_ | ~new_G5185_;
  assign new_G5243_ = ~new_G5239_;
  assign new_G3862_ = ~new_G3860_ | ~new_G3861_;
  assign new_G3871_ = ~new_G3869_ | ~new_G3870_;
  assign new_G3883_ = ~new_G3881_ | ~new_G3882_;
  assign new_G3892_ = ~new_G3890_ | ~new_G3891_;
  assign new_G3956_ = ~new_G3954_ & ~new_G3955_;
  assign new_G3959_ = ~new_G3957_ & ~new_G3958_;
  assign new_G4756_ = new_G1837_ | new_G1875_;
  assign new_G5150_ = ~new_G5145_ | ~new_G5148_;
  assign new_G5151_ = ~new_G5142_ | ~new_G5149_;
  assign new_G5160_ = ~new_G5155_ | ~new_G5158_;
  assign new_G5161_ = ~new_G5152_ | ~new_G5159_;
  assign new_G5194_ = ~new_G5189_ | ~new_G5192_;
  assign new_G5195_ = ~new_G5186_ | ~new_G5193_;
  assign new_G5204_ = ~new_G5199_ | ~new_G5202_;
  assign new_G5205_ = ~new_G5196_ | ~new_G5203_;
  assign new_G5236_ = ~new_G3518_ | ~new_G3515_;
  assign new_G5286_ = new_G3350_;
  assign new_G5379_ = ~new_G5284_ | ~new_G5285_;
  assign new_G5389_ = ~new_G5320_ | ~new_G5321_;
  assign new_G5425_ = ~new_G5404_ | ~new_G5405_;
  assign G610 = new_G609_ & new_G607_ & new_G608_;
  assign new_G1023_ = ~new_G1021_ | ~new_G1022_;
  assign new_G1034_ = ~new_G1032_ | ~new_G1033_;
  assign new_G1052_ = ~new_G1050_ | ~new_G1051_;
  assign new_G1080_ = ~new_G1078_ | ~new_G1079_;
  assign new_G1089_ = ~new_G1087_ | ~new_G1088_;
  assign new_G1100_ = ~new_G1098_ | ~new_G1099_;
  assign new_G1116_ = ~new_G1114_ | ~new_G1115_;
  assign new_G1134_ = ~new_G1132_ | ~new_G1133_;
  assign new_G1152_ = ~new_G1150_ | ~new_G1151_;
  assign new_G4242_ = ~new_G4236_;
  assign new_G1278_ = ~new_G1276_ | ~new_G1277_;
  assign new_G1289_ = ~new_G1287_ | ~new_G1288_;
  assign new_G1307_ = ~new_G1305_ | ~new_G1306_;
  assign new_G1332_ = ~new_G1330_ | ~new_G1331_;
  assign new_G1344_ = ~new_G1342_ | ~new_G1343_;
  assign new_G1365_ = ~new_G1363_ | ~new_G1364_;
  assign new_G1390_ = ~new_G1388_ | ~new_G1389_;
  assign new_G1422_ = ~new_G1420_ | ~new_G1421_;
  assign new_G1430_ = ~new_G1428_ | ~new_G1429_;
  assign new_G1730_ = ~new_G1728_ | ~new_G1729_;
  assign new_G1758_ = ~new_G1756_ | ~new_G1757_;
  assign new_G1767_ = ~new_G1765_ | ~new_G1766_;
  assign new_G1794_ = ~new_G1792_ | ~new_G1793_;
  assign new_G1812_ = ~new_G1810_ | ~new_G1811_;
  assign new_G1876_ = ~new_G4679_ | ~new_G4682_;
  assign new_G4683_ = ~new_G4679_;
  assign new_G4691_ = ~new_G4687_;
  assign new_G4699_ = ~new_G4695_;
  assign new_G4707_ = ~new_G4703_;
  assign new_G4715_ = ~new_G4711_;
  assign new_G4730_ = ~new_G4724_;
  assign new_G1984_ = ~new_G1982_ | ~new_G1983_;
  assign new_G2009_ = ~new_G2007_ | ~new_G2008_;
  assign new_G2042_ = ~new_G2040_ | ~new_G2041_;
  assign new_G2067_ = ~new_G2065_ | ~new_G2066_;
  assign new_G2099_ = ~new_G2097_ | ~new_G2098_;
  assign new_G4869_ = ~new_G4865_;
  assign new_G4927_ = ~new_G4923_;
  assign new_G3445_ = ~new_G3443_ | ~new_G3444_;
  assign new_G3454_ = ~new_G3452_ | ~new_G3453_;
  assign new_G3463_ = ~new_G3461_ | ~new_G3462_;
  assign new_G3468_ = ~new_G3466_ | ~new_G3467_;
  assign new_G3477_ = ~new_G3475_ | ~new_G3476_;
  assign new_G3486_ = ~new_G3484_ | ~new_G3485_;
  assign new_G4103_ = new_G4099_ & new_G3170_;
  assign new_G4412_ = ~new_G4406_;
  assign new_G4558_ = ~new_G4552_;
  assign new_G4859_ = ~new_G4855_;
  assign new_G4876_ = ~new_G4870_;
  assign new_G4917_ = ~new_G4913_;
  assign new_G4955_ = ~new_G4951_;
  assign new_G5012_ = ~new_G5006_;
  assign new_G5043_ = ~new_G5039_;
  assign new_G5216_ = ~new_G5160_ | ~new_G5161_;
  assign new_G5219_ = ~new_G5150_ | ~new_G5151_;
  assign new_G5226_ = ~new_G5204_ | ~new_G5205_;
  assign new_G5229_ = ~new_G5194_ | ~new_G5195_;
  assign new_G5392_ = ~new_G5386_;
  assign new_G5422_ = ~new_G3959_ | ~new_G3956_;
  assign new_G1866_ = new_G1778_ & new_G1806_;
  assign new_G1877_ = ~new_G4676_ | ~new_G4683_;
  assign new_G4762_ = ~new_G4756_;
  assign new_G2142_ = new_G2021_ & new_G2059_;
  assign new_G2146_ = new_G2021_ & new_G2059_;
  assign new_G5242_ = ~new_G5236_;
  assign new_G3532_ = ~new_G5236_ | ~new_G5243_;
  assign new_G3866_ = ~new_G3862_;
  assign new_G3887_ = ~new_G3883_;
  assign new_G3918_ = new_G3871_;
  assign new_G3922_ = new_G3871_;
  assign new_G3926_ = new_G3892_;
  assign new_G3930_ = new_G3892_;
  assign new_G5429_ = ~new_G5425_;
  assign new_G4104_ = new_G4099_ | new_G4103_;
  assign new_G4743_ = new_G1778_;
  assign new_G4991_ = new_G2021_;
  assign new_G5001_ = new_G2021_;
  assign new_G5292_ = ~new_G5286_;
  assign new_G5295_ = ~new_G5286_ | ~new_G5293_;
  assign new_G5383_ = ~new_G5379_;
  assign new_G5393_ = ~new_G5389_;
  assign new_G5394_ = ~new_G5389_ | ~new_G5392_;
  assign new_G1439_ = new_G1278_ & new_G1301_;
  assign new_G1440_ = new_G1318_ & new_G1289_ & new_G1278_;
  assign new_G1441_ = new_G1289_ & new_G1324_ & new_G1307_ & new_G1278_;
  assign new_G1847_ = new_G1712_ & new_G1749_ & new_G1730_ & new_G1704_;
  assign new_G1168_ = new_G1023_ & new_G1046_;
  assign new_G1169_ = new_G1064_ & new_G1034_ & new_G1023_;
  assign new_G1170_ = new_G1034_ & new_G1071_ & new_G1052_ & new_G1023_;
  assign new_G2117_ = new_G1966_ & new_G2001_ & new_G1984_ & new_G1958_;
  assign new_G1086_ = ~new_G1080_;
  assign new_G1166_ = new_G1023_ & new_G1052_ & new_G1034_ & new_G1080_;
  assign new_G1171_ = new_G1034_ & new_G1064_;
  assign new_G1172_ = new_G1034_ & new_G1052_ & new_G1071_;
  assign new_G1173_ = new_G1034_ & new_G1080_ & new_G1052_;
  assign new_G1174_ = new_G1034_ & new_G1064_;
  assign new_G1175_ = new_G1034_ & new_G1071_ & new_G1052_;
  assign new_G1176_ = new_G1052_ & new_G1071_;
  assign new_G1177_ = new_G1080_ & new_G1052_;
  assign new_G1178_ = new_G1052_ & new_G1071_;
  assign new_G1179_ = new_G1134_ & new_G1089_ & new_G1116_ & new_G1100_ & new_G1152_;
  assign new_G1181_ = new_G1089_ & new_G1111_;
  assign new_G1182_ = new_G1128_ & new_G1100_ & new_G1089_;
  assign new_G1183_ = new_G1100_ & new_G1145_ & new_G1116_ & new_G1089_;
  assign new_G1184_ = new_G1100_ & new_G1160_ & new_G1089_ & new_G1134_ & new_G1116_;
  assign new_G1188_ = new_G1100_ & new_G1128_;
  assign new_G1189_ = new_G1100_ & new_G1116_ & new_G1145_;
  assign new_G1190_ = new_G1100_ & new_G1160_ & new_G1134_ & new_G1116_;
  assign new_G1191_ = new_G1100_ & new_G1134_ & new_G1116_ & G4 & new_G1152_;
  assign new_G1192_ = new_G1145_ & new_G1116_;
  assign new_G1193_ = new_G1160_ & new_G1134_ & new_G1116_;
  assign new_G1194_ = new_G1134_ & new_G1116_ & G4 & new_G1152_;
  assign new_G1195_ = new_G1134_ & new_G1160_;
  assign new_G1196_ = new_G1134_ & G4 & new_G1152_;
  assign new_G1197_ = G4 & new_G1152_;
  assign new_G1437_ = new_G1278_ & new_G1289_ & new_G1422_ & new_G1307_;
  assign new_G1442_ = new_G1289_ & new_G1318_;
  assign new_G1443_ = new_G1289_ & new_G1307_ & new_G1324_;
  assign new_G1444_ = new_G1289_ & new_G1422_ & new_G1307_;
  assign new_G1445_ = new_G1289_ & new_G1318_;
  assign new_G1446_ = new_G1289_ & new_G1307_ & new_G1324_;
  assign new_G1447_ = new_G1307_ & new_G1324_;
  assign new_G1451_ = new_G1332_ & new_G1344_ & new_G1365_ & new_G1430_ & new_G1390_;
  assign new_G1454_ = new_G1332_ & new_G1359_;
  assign new_G1455_ = new_G1382_ & new_G1344_ & new_G1332_;
  assign new_G1456_ = new_G1344_ & new_G1404_ & new_G1365_ & new_G1332_;
  assign new_G1457_ = new_G1344_ & new_G1412_ & new_G1332_ & new_G1390_ & new_G1365_;
  assign new_G1465_ = new_G1344_ & new_G1382_;
  assign new_G1466_ = new_G1344_ & new_G1365_ & new_G1404_;
  assign new_G1467_ = new_G1344_ & new_G1412_ & new_G1390_ & new_G1365_;
  assign new_G1468_ = new_G1390_ & new_G1344_ & new_G1430_ & new_G1365_;
  assign new_G1469_ = new_G1344_ & new_G1382_;
  assign new_G1470_ = new_G1344_ & new_G1365_ & new_G1404_;
  assign new_G1471_ = new_G1344_ & new_G1412_ & new_G1390_ & new_G1365_;
  assign new_G1472_ = new_G1365_ & new_G1404_;
  assign new_G1473_ = new_G1412_ & new_G1390_ & new_G1365_;
  assign new_G1474_ = new_G1390_ & new_G1430_ & new_G1365_;
  assign new_G1475_ = new_G1365_ & new_G1404_;
  assign new_G1476_ = new_G1412_ & new_G1390_ & new_G1365_;
  assign new_G1477_ = new_G1390_ & new_G1412_;
  assign new_G1481_ = new_G1422_ & new_G1307_;
  assign new_G1482_ = new_G1430_ & new_G1390_;
  assign new_G1764_ = ~new_G1758_;
  assign new_G1843_ = new_G1704_ & new_G1730_ & new_G1712_ & new_G1758_;
  assign new_G1850_ = new_G1712_ & new_G1730_ & new_G1749_;
  assign new_G1851_ = new_G1712_ & new_G1758_ & new_G1730_;
  assign new_G1853_ = new_G1712_ & new_G1749_ & new_G1730_;
  assign new_G1854_ = new_G1730_ & new_G1749_;
  assign new_G1855_ = new_G1758_ & new_G1730_;
  assign new_G1856_ = new_G1730_ & new_G1749_;
  assign new_G1857_ = new_G1812_ & new_G1767_ & new_G1794_ & new_G1778_ & new_G1829_;
  assign new_G1859_ = new_G1767_ & new_G1789_;
  assign new_G1860_ = new_G1806_ & new_G1778_ & new_G1767_;
  assign new_G1861_ = new_G1778_ & new_G1823_ & new_G1794_ & new_G1767_;
  assign new_G1862_ = new_G1778_ & new_G1837_ & new_G1767_ & new_G1812_ & new_G1794_;
  assign new_G1867_ = new_G1778_ & new_G1794_ & new_G1823_;
  assign new_G1868_ = new_G1778_ & new_G1837_ & new_G1812_ & new_G1794_;
  assign new_G1869_ = new_G1778_ & new_G1812_ & new_G1794_ & G54 & new_G1829_;
  assign new_G1870_ = new_G1823_ & new_G1794_;
  assign new_G1871_ = new_G1837_ & new_G1812_ & new_G1794_;
  assign new_G1872_ = new_G1812_ & new_G1794_ & G54 & new_G1829_;
  assign new_G1873_ = new_G1812_ & new_G1837_;
  assign new_G1874_ = new_G1812_ & G54 & new_G1829_;
  assign new_G1878_ = ~new_G1876_ | ~new_G1877_;
  assign new_G2113_ = new_G1958_ & new_G1966_ & new_G2099_ & new_G1984_;
  assign new_G2120_ = new_G1966_ & new_G1984_ & new_G2001_;
  assign new_G2121_ = new_G1966_ & new_G2099_ & new_G1984_;
  assign new_G2123_ = new_G1966_ & new_G1984_ & new_G2001_;
  assign new_G2124_ = new_G1984_ & new_G2001_;
  assign new_G2128_ = new_G2009_ & new_G2021_ & new_G2042_ & new_G2106_ & new_G2067_;
  assign new_G2131_ = new_G2009_ & new_G2036_;
  assign new_G2132_ = new_G2059_ & new_G2021_ & new_G2009_;
  assign new_G2133_ = new_G2021_ & new_G2081_ & new_G2042_ & new_G2009_;
  assign new_G2134_ = new_G2021_ & new_G2089_ & new_G2009_ & new_G2067_ & new_G2042_;
  assign new_G2143_ = new_G2021_ & new_G2042_ & new_G2081_;
  assign new_G2144_ = new_G2021_ & new_G2089_ & new_G2067_ & new_G2042_;
  assign new_G2145_ = new_G2067_ & new_G2021_ & new_G2106_ & new_G2042_;
  assign new_G2147_ = new_G2021_ & new_G2042_ & new_G2081_;
  assign new_G2148_ = new_G2021_ & new_G2089_ & new_G2067_ & new_G2042_;
  assign new_G2149_ = new_G2042_ & new_G2081_;
  assign new_G2150_ = new_G2089_ & new_G2067_ & new_G2042_;
  assign new_G2151_ = new_G2067_ & new_G2106_ & new_G2042_;
  assign new_G2152_ = new_G2042_ & new_G2081_;
  assign new_G2153_ = new_G2089_ & new_G2067_ & new_G2042_;
  assign new_G2154_ = new_G2067_ & new_G2089_;
  assign new_G2158_ = new_G2099_ & new_G1984_;
  assign new_G2159_ = new_G2106_ & new_G2067_;
  assign new_G3449_ = ~new_G3445_;
  assign new_G3458_ = ~new_G3454_;
  assign new_G3472_ = ~new_G3468_;
  assign new_G3481_ = ~new_G3477_;
  assign new_G3497_ = new_G3463_;
  assign new_G3501_ = new_G3463_;
  assign new_G3505_ = new_G3486_;
  assign new_G3509_ = new_G3486_;
  assign new_G3531_ = ~new_G5239_ | ~new_G5242_;
  assign new_G5428_ = ~new_G5422_;
  assign new_G3967_ = ~new_G5422_ | ~new_G5429_;
  assign new_G4191_ = new_G1152_;
  assign new_G4199_ = new_G1023_;
  assign new_G4207_ = new_G1023_;
  assign new_G4215_ = new_G1034_;
  assign new_G4223_ = new_G1034_;
  assign new_G4231_ = new_G1052_;
  assign new_G4239_ = new_G1052_;
  assign new_G4247_ = new_G1089_;
  assign new_G4255_ = new_G1100_;
  assign new_G4263_ = new_G1116_;
  assign new_G4271_ = new_G1134_;
  assign new_G4371_ = new_G1422_;
  assign new_G4381_ = new_G1307_;
  assign new_G4391_ = new_G1278_;
  assign new_G4401_ = new_G1289_;
  assign new_G4429_ = new_G1422_;
  assign new_G4439_ = new_G1307_;
  assign new_G4449_ = new_G1278_;
  assign new_G4459_ = new_G1289_;
  assign new_G4497_ = new_G1430_;
  assign new_G4507_ = new_G1390_;
  assign new_G4517_ = new_G1332_;
  assign new_G4527_ = new_G1365_;
  assign new_G4537_ = new_G1344_;
  assign new_G4547_ = new_G1344_;
  assign new_G4585_ = new_G1430_;
  assign new_G4595_ = new_G1390_;
  assign new_G4605_ = new_G1332_;
  assign new_G4615_ = new_G1365_;
  assign new_G4719_ = new_G1730_;
  assign new_G4727_ = new_G1730_;
  assign new_G4735_ = new_G1767_;
  assign new_G4751_ = new_G1794_;
  assign new_G4759_ = new_G1812_;
  assign new_G4835_ = new_G2099_;
  assign new_G4845_ = new_G1984_;
  assign new_G4893_ = new_G2099_;
  assign new_G4903_ = new_G1984_;
  assign new_G4961_ = new_G2067_;
  assign new_G4971_ = new_G2009_;
  assign new_G4981_ = new_G2042_;
  assign new_G5049_ = new_G2067_;
  assign new_G5059_ = new_G2009_;
  assign new_G5069_ = new_G2042_;
  assign new_G5222_ = ~new_G5216_;
  assign new_G5223_ = ~new_G5219_;
  assign new_G5232_ = ~new_G5226_;
  assign new_G5233_ = ~new_G5229_;
  assign new_G5294_ = ~new_G5289_ | ~new_G5292_;
  assign new_G5395_ = ~new_G5386_ | ~new_G5393_;
  assign new_G589_ = new_G1441_ | new_G1440_ | new_G1286_ | new_G1439_;
  assign new_G616_ = new_G1847_ | new_G1846_ | new_G3167_ | new_G1845_;
  assign new_G619_ = new_G1170_ | new_G1169_ | new_G1031_ | new_G1168_;
  assign new_G627_ = new_G2117_ | new_G2116_ | new_G3167_ | new_G2115_;
  assign new_G1185_ = new_G1184_ | new_G1183_ | new_G1182_ | new_G1097_ | new_G1181_;
  assign new_G1448_ = new_G1318_ | new_G1447_;
  assign new_G1458_ = new_G1457_ | new_G1456_ | new_G1455_ | new_G1341_ | new_G1454_;
  assign new_G1478_ = new_G1404_ | new_G1477_;
  assign new_G1863_ = new_G1862_ | new_G1861_ | new_G1860_ | new_G1775_ | new_G1859_;
  assign new_G4747_ = ~new_G4743_;
  assign new_G2125_ = new_G1995_ | new_G2124_;
  assign new_G2135_ = new_G2134_ | new_G2133_ | new_G2132_ | new_G2018_ | new_G2131_;
  assign new_G2155_ = new_G2081_ | new_G2154_;
  assign new_G4995_ = ~new_G4991_;
  assign new_G5005_ = ~new_G5001_;
  assign new_G3533_ = ~new_G3531_ | ~new_G3532_;
  assign new_G3921_ = ~new_G3918_;
  assign new_G3925_ = ~new_G3922_;
  assign new_G3929_ = ~new_G3926_;
  assign new_G3933_ = ~new_G3930_;
  assign new_G3943_ = new_G3918_ & new_G3862_ & new_G3853_;
  assign new_G3946_ = new_G3922_ & new_G3866_ & new_G3857_;
  assign new_G3949_ = new_G3926_ & new_G3883_ & new_G3874_;
  assign new_G3952_ = new_G3930_ & new_G3887_ & new_G3878_;
  assign new_G3966_ = ~new_G5425_ | ~new_G5428_;
  assign new_G4107_ = ~new_G4104_ | ~G132;
  assign new_G4196_ = new_G1173_ | new_G1172_ | new_G1046_ | new_G1171_;
  assign new_G4204_ = ~new_G1175_ & ~new_G1046_ & ~new_G1174_;
  assign new_G4212_ = new_G1177_ | new_G1064_ | new_G1176_;
  assign new_G4220_ = ~new_G1064_ & ~new_G1178_;
  assign new_G4244_ = new_G1191_ | new_G1190_ | new_G1189_ | new_G1111_ | new_G1188_;
  assign new_G4252_ = new_G1194_ | new_G1193_ | new_G1128_ | new_G1192_;
  assign new_G4260_ = new_G1196_ | new_G1145_ | new_G1195_;
  assign new_G4268_ = new_G1160_ | new_G1197_;
  assign new_G4361_ = new_G1444_ | new_G1443_ | new_G1301_ | new_G1442_;
  assign new_G4419_ = ~new_G1446_ & ~new_G1301_ & ~new_G1445_;
  assign new_G4467_ = new_G1474_ | new_G1473_ | new_G1382_ | new_G1472_;
  assign new_G4487_ = new_G1468_ | new_G1467_ | new_G1466_ | new_G1359_ | new_G1465_;
  assign new_G4555_ = ~new_G1476_ & ~new_G1382_ & ~new_G1475_;
  assign new_G4575_ = ~new_G1471_ & ~new_G1470_ & ~new_G1359_ & ~new_G1469_;
  assign new_G4684_ = new_G1851_ | new_G1850_ | new_G1724_ | new_G1849_;
  assign new_G4692_ = ~new_G1853_ & ~new_G1724_ & ~new_G1852_;
  assign new_G4700_ = new_G1855_ | new_G1742_ | new_G1854_;
  assign new_G4708_ = ~new_G1742_ & ~new_G1856_;
  assign new_G4732_ = new_G1869_ | new_G1868_ | new_G1867_ | new_G1789_ | new_G1866_;
  assign new_G4740_ = new_G1872_ | new_G1871_ | new_G1806_ | new_G1870_;
  assign new_G4748_ = new_G1874_ | new_G1823_ | new_G1873_;
  assign new_G4825_ = new_G2121_ | new_G2120_ | new_G1978_ | new_G2119_;
  assign new_G4883_ = ~new_G2123_ & ~new_G1978_ & ~new_G2122_;
  assign new_G4928_ = new_G2151_ | new_G2150_ | new_G2059_ | new_G2149_;
  assign new_G4941_ = new_G2145_ | new_G2144_ | new_G2143_ | new_G2036_ | new_G2142_;
  assign new_G5009_ = ~new_G2153_ & ~new_G2059_ & ~new_G2152_;
  assign new_G5029_ = ~new_G2148_ & ~new_G2147_ & ~new_G2036_ & ~new_G2146_;
  assign new_G5224_ = ~new_G5219_ | ~new_G5222_;
  assign new_G5225_ = ~new_G5216_ | ~new_G5223_;
  assign new_G5234_ = ~new_G5229_ | ~new_G5232_;
  assign new_G5235_ = ~new_G5226_ | ~new_G5233_;
  assign new_G5376_ = ~new_G5294_ | ~new_G5295_;
  assign new_G5417_ = ~new_G5394_ | ~new_G5395_;
  assign new_G576_ = ~new_G1878_;
  assign G588 = new_G1437_ & new_G1451_;
  assign G615 = new_G1843_ & new_G1857_;
  assign G626 = new_G2113_ & new_G2128_;
  assign G632 = new_G1166_ & new_G1179_;
  assign new_G1198_ = ~new_G4191_ | ~new_G4194_;
  assign new_G4195_ = ~new_G4191_;
  assign new_G4203_ = ~new_G4199_;
  assign new_G4211_ = ~new_G4207_;
  assign new_G4219_ = ~new_G4215_;
  assign new_G4227_ = ~new_G4223_;
  assign new_G1217_ = ~new_G4231_ | ~new_G4234_;
  assign new_G4235_ = ~new_G4231_;
  assign new_G1221_ = ~new_G4239_ | ~new_G4242_;
  assign new_G4243_ = ~new_G4239_;
  assign new_G1224_ = new_G1179_ & G4;
  assign new_G4251_ = ~new_G4247_;
  assign new_G4259_ = ~new_G4255_;
  assign new_G4267_ = ~new_G4263_;
  assign new_G4275_ = ~new_G4271_;
  assign new_G1453_ = ~new_G1451_;
  assign new_G4405_ = ~new_G4401_;
  assign new_G4463_ = ~new_G4459_;
  assign new_G4541_ = ~new_G4537_;
  assign new_G4551_ = ~new_G4547_;
  assign new_G1895_ = ~new_G4719_ | ~new_G4722_;
  assign new_G4723_ = ~new_G4719_;
  assign new_G1899_ = ~new_G4727_ | ~new_G4730_;
  assign new_G4731_ = ~new_G4727_;
  assign new_G1902_ = new_G1857_ & G54;
  assign new_G4739_ = ~new_G4735_;
  assign new_G4755_ = ~new_G4751_;
  assign new_G1929_ = ~new_G4759_ | ~new_G4762_;
  assign new_G4763_ = ~new_G4759_;
  assign new_G2130_ = ~new_G2128_;
  assign new_G3500_ = ~new_G3497_;
  assign new_G3504_ = ~new_G3501_;
  assign new_G3508_ = ~new_G3505_;
  assign new_G3512_ = ~new_G3509_;
  assign new_G3520_ = new_G3497_ & new_G3454_ & new_G3445_;
  assign new_G3523_ = new_G3501_ & new_G3458_ & new_G3449_;
  assign new_G3526_ = new_G3505_ & new_G3477_ & new_G3468_;
  assign new_G3529_ = new_G3509_ & new_G3481_ & new_G3472_;
  assign G1002 = new_G3533_;
  assign new_G3837_ = new_G3823_ & new_G1878_ & new_G3795_;
  assign new_G3942_ = new_G3921_ & new_G3857_ & new_G3862_;
  assign new_G3945_ = new_G3925_ & new_G3853_ & new_G3866_;
  assign new_G3948_ = new_G3929_ & new_G3878_ & new_G3883_;
  assign new_G3951_ = new_G3933_ & new_G3874_ & new_G3887_;
  assign new_G3968_ = ~new_G3966_ | ~new_G3967_;
  assign new_G4375_ = ~new_G4371_;
  assign new_G4385_ = ~new_G4381_;
  assign new_G4395_ = ~new_G4391_;
  assign new_G4433_ = ~new_G4429_;
  assign new_G4443_ = ~new_G4439_;
  assign new_G4453_ = ~new_G4449_;
  assign new_G4501_ = ~new_G4497_;
  assign new_G4511_ = ~new_G4507_;
  assign new_G4521_ = ~new_G4517_;
  assign new_G4531_ = ~new_G4527_;
  assign new_G4619_ = ~new_G4615_;
  assign new_G4589_ = ~new_G4585_;
  assign new_G4599_ = ~new_G4595_;
  assign new_G4609_ = ~new_G4605_;
  assign new_G4839_ = ~new_G4835_;
  assign new_G4849_ = ~new_G4845_;
  assign new_G4897_ = ~new_G4893_;
  assign new_G4907_ = ~new_G4903_;
  assign new_G4965_ = ~new_G4961_;
  assign new_G4975_ = ~new_G4971_;
  assign new_G4985_ = ~new_G4981_;
  assign new_G5073_ = ~new_G5069_;
  assign new_G5053_ = ~new_G5049_;
  assign new_G5063_ = ~new_G5059_;
  assign new_G5247_ = ~new_G5224_ | ~new_G5225_;
  assign new_G5255_ = ~new_G5234_ | ~new_G5235_;
  assign new_G590_ = new_G1437_ & new_G1458_;
  assign new_G617_ = new_G1863_ & new_G1843_;
  assign new_G620_ = new_G1185_ & new_G1166_;
  assign new_G628_ = new_G2113_ & new_G2135_;
  assign new_G3535_ = ~new_G3533_;
  assign new_G1199_ = ~new_G4188_ | ~new_G4195_;
  assign new_G4202_ = ~new_G4196_;
  assign new_G1204_ = ~new_G4196_ | ~new_G4203_;
  assign new_G4210_ = ~new_G4204_;
  assign new_G1207_ = ~new_G4204_ | ~new_G4211_;
  assign new_G4218_ = ~new_G4212_;
  assign new_G1211_ = ~new_G4212_ | ~new_G4219_;
  assign new_G4226_ = ~new_G4220_;
  assign new_G1214_ = ~new_G4220_ | ~new_G4227_;
  assign new_G1218_ = ~new_G4228_ | ~new_G4235_;
  assign new_G1222_ = ~new_G4236_ | ~new_G4243_;
  assign new_G1225_ = new_G1185_ | new_G1224_;
  assign new_G4250_ = ~new_G4244_;
  assign new_G1237_ = ~new_G4244_ | ~new_G4251_;
  assign new_G4258_ = ~new_G4252_;
  assign new_G1242_ = ~new_G4252_ | ~new_G4259_;
  assign new_G4266_ = ~new_G4260_;
  assign new_G1247_ = ~new_G4260_ | ~new_G4267_;
  assign new_G4274_ = ~new_G4268_;
  assign new_G1252_ = ~new_G4268_ | ~new_G4275_;
  assign new_G1462_ = ~new_G1458_;
  assign new_G4690_ = ~new_G4684_;
  assign new_G1882_ = ~new_G4684_ | ~new_G4691_;
  assign new_G4698_ = ~new_G4692_;
  assign new_G1885_ = ~new_G4692_ | ~new_G4699_;
  assign new_G4706_ = ~new_G4700_;
  assign new_G1889_ = ~new_G4700_ | ~new_G4707_;
  assign new_G4714_ = ~new_G4708_;
  assign new_G1892_ = ~new_G4708_ | ~new_G4715_;
  assign new_G1896_ = ~new_G4716_ | ~new_G4723_;
  assign new_G1900_ = ~new_G4724_ | ~new_G4731_;
  assign new_G1903_ = new_G1863_ | new_G1902_;
  assign new_G4738_ = ~new_G4732_;
  assign new_G1915_ = ~new_G4732_ | ~new_G4739_;
  assign new_G4746_ = ~new_G4740_;
  assign new_G1920_ = ~new_G4740_ | ~new_G4747_;
  assign new_G4754_ = ~new_G4748_;
  assign new_G1925_ = ~new_G4748_ | ~new_G4755_;
  assign new_G1930_ = ~new_G4756_ | ~new_G4763_;
  assign new_G2139_ = ~new_G2135_;
  assign new_G3519_ = new_G3500_ & new_G3449_ & new_G3454_;
  assign new_G3522_ = new_G3504_ & new_G3445_ & new_G3458_;
  assign new_G3525_ = new_G3508_ & new_G3472_ & new_G3477_;
  assign new_G3528_ = new_G3512_ & new_G3468_ & new_G3481_;
  assign new_G3848_ = new_G3838_ | new_G3836_ | new_G3837_;
  assign new_G3944_ = ~new_G3942_ & ~new_G3943_;
  assign new_G3947_ = ~new_G3945_ & ~new_G3946_;
  assign new_G3950_ = ~new_G3948_ & ~new_G3949_;
  assign new_G3953_ = ~new_G3951_ & ~new_G3952_;
  assign new_G5421_ = ~new_G5417_;
  assign G1004 = new_G3968_;
  assign new_G4111_ = new_G4104_ & new_G4107_;
  assign new_G4112_ = new_G4107_ & G132;
  assign new_G4351_ = new_G1448_ | new_G1481_;
  assign new_G4365_ = ~new_G4361_;
  assign new_G4409_ = ~new_G1448_;
  assign new_G4423_ = ~new_G4419_;
  assign new_G4471_ = ~new_G4467_;
  assign new_G4472_ = ~new_G4467_ | ~new_G4470_;
  assign new_G4477_ = new_G1478_ | new_G1482_;
  assign new_G4491_ = ~new_G4487_;
  assign new_G4559_ = ~new_G4555_;
  assign new_G4560_ = ~new_G4555_ | ~new_G4558_;
  assign new_G4565_ = ~new_G1478_;
  assign new_G4579_ = ~new_G4575_;
  assign new_G4815_ = new_G2125_ | new_G2158_;
  assign new_G4829_ = ~new_G4825_;
  assign new_G4873_ = ~new_G2125_;
  assign new_G4887_ = ~new_G4883_;
  assign new_G4931_ = new_G2155_ | new_G2159_;
  assign new_G4934_ = ~new_G4928_;
  assign new_G4945_ = ~new_G4941_;
  assign new_G5013_ = ~new_G5009_;
  assign new_G5014_ = ~new_G5009_ | ~new_G5012_;
  assign new_G5019_ = ~new_G2155_;
  assign new_G5033_ = ~new_G5029_;
  assign new_G5382_ = ~new_G5376_;
  assign new_G5385_ = ~new_G5376_ | ~new_G5383_;
  assign G591 = new_G589_ | new_G590_;
  assign G618 = new_G616_ | new_G617_;
  assign G621 = new_G619_ | new_G620_;
  assign G629 = new_G627_ | new_G628_;
  assign new_G3970_ = ~new_G3968_;
  assign new_G1200_ = ~new_G1198_ | ~new_G1199_;
  assign new_G1203_ = ~new_G4199_ | ~new_G4202_;
  assign new_G1206_ = ~new_G4207_ | ~new_G4210_;
  assign new_G1210_ = ~new_G4215_ | ~new_G4218_;
  assign new_G1213_ = ~new_G4223_ | ~new_G4226_;
  assign new_G1219_ = ~new_G1217_ | ~new_G1218_;
  assign new_G1223_ = ~new_G1221_ | ~new_G1222_;
  assign new_G1236_ = ~new_G4247_ | ~new_G4250_;
  assign new_G1241_ = ~new_G4255_ | ~new_G4258_;
  assign new_G1246_ = ~new_G4263_ | ~new_G4266_;
  assign new_G1251_ = ~new_G4271_ | ~new_G4274_;
  assign new_G1881_ = ~new_G4687_ | ~new_G4690_;
  assign new_G1884_ = ~new_G4695_ | ~new_G4698_;
  assign new_G1888_ = ~new_G4703_ | ~new_G4706_;
  assign new_G1891_ = ~new_G4711_ | ~new_G4714_;
  assign new_G1897_ = ~new_G1895_ | ~new_G1896_;
  assign new_G1901_ = ~new_G1899_ | ~new_G1900_;
  assign new_G1914_ = ~new_G4735_ | ~new_G4738_;
  assign new_G1919_ = ~new_G4743_ | ~new_G4746_;
  assign new_G1924_ = ~new_G4751_ | ~new_G4754_;
  assign new_G1931_ = ~new_G1929_ | ~new_G1930_;
  assign new_G3521_ = ~new_G3519_ & ~new_G3520_;
  assign new_G3524_ = ~new_G3522_ & ~new_G3523_;
  assign new_G3527_ = ~new_G3525_ & ~new_G3526_;
  assign new_G3530_ = ~new_G3528_ & ~new_G3529_;
  assign new_G5251_ = ~new_G5247_;
  assign new_G5259_ = ~new_G5255_;
  assign new_G4113_ = new_G4111_ | new_G4112_;
  assign new_G4473_ = ~new_G4464_ | ~new_G4471_;
  assign new_G4561_ = ~new_G4552_ | ~new_G4559_;
  assign new_G5015_ = ~new_G5006_ | ~new_G5013_;
  assign new_G5384_ = ~new_G5379_ | ~new_G5382_;
  assign new_G5406_ = ~new_G3947_ | ~new_G3944_;
  assign new_G5414_ = ~new_G3953_ | ~new_G3950_;
  assign new_G1664_ = new_G1645_ & new_G3848_ & new_G1621_;
  assign new_G2335_ = new_G2316_ & new_G3848_ & new_G2293_;
  assign new_G718_ = new_G2454_ & new_G3848_ & new_G2430_;
  assign G822 = ~new_G3848_;
  assign new_G855_ = new_G2512_ & new_G3848_ & new_G2488_;
  assign new_G1205_ = ~new_G1203_ | ~new_G1204_;
  assign new_G1208_ = ~new_G1206_ | ~new_G1207_;
  assign new_G1212_ = ~new_G1210_ | ~new_G1211_;
  assign new_G1215_ = ~new_G1213_ | ~new_G1214_;
  assign new_G1220_ = ~new_G1219_;
  assign new_G1231_ = ~new_G1225_;
  assign new_G1238_ = ~new_G1236_ | ~new_G1237_;
  assign new_G1243_ = ~new_G1241_ | ~new_G1242_;
  assign new_G1248_ = ~new_G1246_ | ~new_G1247_;
  assign new_G1253_ = ~new_G1251_ | ~new_G1252_;
  assign new_G1272_ = new_G1225_ & new_G1086_;
  assign new_G1483_ = new_G1462_ & new_G1453_;
  assign new_G1883_ = ~new_G1881_ | ~new_G1882_;
  assign new_G1886_ = ~new_G1884_ | ~new_G1885_;
  assign new_G1890_ = ~new_G1888_ | ~new_G1889_;
  assign new_G1893_ = ~new_G1891_ | ~new_G1892_;
  assign new_G1898_ = ~new_G1897_;
  assign new_G1909_ = ~new_G1903_;
  assign new_G1916_ = ~new_G1914_ | ~new_G1915_;
  assign new_G1921_ = ~new_G1919_ | ~new_G1920_;
  assign new_G1926_ = ~new_G1924_ | ~new_G1925_;
  assign new_G1953_ = new_G1903_ & new_G1764_;
  assign new_G2160_ = new_G2139_ & new_G2130_;
  assign new_G4355_ = ~new_G4351_;
  assign new_G4356_ = ~new_G4351_ | ~new_G4354_;
  assign new_G4413_ = ~new_G4409_;
  assign new_G4414_ = ~new_G4409_ | ~new_G4412_;
  assign new_G4474_ = ~new_G4472_ | ~new_G4473_;
  assign new_G4481_ = ~new_G4477_;
  assign new_G4562_ = ~new_G4560_ | ~new_G4561_;
  assign new_G4569_ = ~new_G4565_;
  assign new_G4819_ = ~new_G4815_;
  assign new_G4820_ = ~new_G4815_ | ~new_G4818_;
  assign new_G4877_ = ~new_G4873_;
  assign new_G4878_ = ~new_G4873_ | ~new_G4876_;
  assign new_G4935_ = ~new_G4931_;
  assign new_G4936_ = ~new_G4931_ | ~new_G4934_;
  assign new_G5016_ = ~new_G5014_ | ~new_G5015_;
  assign new_G5023_ = ~new_G5019_;
  assign new_G5244_ = ~new_G3524_ | ~new_G3521_;
  assign new_G5252_ = ~new_G3530_ | ~new_G3527_;
  assign new_G5409_ = ~new_G5384_ | ~new_G5385_;
  assign new_G566_ = ~new_G1200_;
  assign new_G577_ = ~new_G1931_;
  assign new_G3733_ = new_G3721_ & new_G4113_ & G3724;
  assign new_G1209_ = ~new_G1208_;
  assign new_G1216_ = ~new_G1215_;
  assign new_G1257_ = new_G1225_ & new_G1205_;
  assign new_G1262_ = new_G1225_ & new_G1212_;
  assign new_G1267_ = new_G1225_ & new_G1220_;
  assign new_G1887_ = ~new_G1886_;
  assign new_G1894_ = ~new_G1893_;
  assign new_G1935_ = new_G1903_ & new_G1883_;
  assign new_G1943_ = new_G1903_ & new_G1890_;
  assign new_G1948_ = new_G1903_ & new_G1898_;
  assign new_G3779_ = new_G3765_ & new_G1200_ & new_G3737_;
  assign new_G3840_ = new_G3823_ & new_G1931_ & new_G3795_;
  assign new_G5412_ = ~new_G5406_;
  assign new_G5420_ = ~new_G5414_;
  assign new_G3964_ = ~new_G5414_ | ~new_G5421_;
  assign new_G4357_ = ~new_G4348_ | ~new_G4355_;
  assign new_G4415_ = ~new_G4406_ | ~new_G4413_;
  assign new_G4821_ = ~new_G4812_ | ~new_G4819_;
  assign new_G4879_ = ~new_G4870_ | ~new_G4877_;
  assign new_G4937_ = ~new_G4928_ | ~new_G4935_;
  assign new_G567_ = ~new_G1253_;
  assign new_G568_ = ~new_G1248_;
  assign new_G569_ = ~new_G1243_;
  assign new_G570_ = ~new_G1238_;
  assign new_G578_ = ~new_G1926_;
  assign new_G579_ = ~new_G1921_;
  assign new_G580_ = ~new_G1916_;
  assign new_G1256_ = new_G1209_ & new_G1231_;
  assign new_G1261_ = new_G1216_ & new_G1231_;
  assign new_G1266_ = new_G1223_ & new_G1231_;
  assign new_G1271_ = new_G1080_ & new_G1231_;
  assign new_G1486_ = ~new_G1483_;
  assign new_G1934_ = new_G1887_ & new_G1909_;
  assign new_G1942_ = new_G1894_ & new_G1909_;
  assign new_G1947_ = new_G1901_ & new_G1909_;
  assign new_G1952_ = new_G1758_ & new_G1909_;
  assign new_G2163_ = ~new_G2160_;
  assign new_G5250_ = ~new_G5244_;
  assign new_G3537_ = ~new_G5244_ | ~new_G5251_;
  assign new_G5258_ = ~new_G5252_;
  assign new_G3542_ = ~new_G5252_ | ~new_G5259_;
  assign new_G3782_ = new_G3765_ & new_G1253_ & new_G3737_;
  assign new_G3785_ = new_G3765_ & new_G1248_ & new_G3737_;
  assign new_G3788_ = new_G3765_ & new_G1243_ & new_G3737_;
  assign new_G3790_ = new_G3780_ | new_G3778_ | new_G3779_;
  assign new_G3843_ = new_G3823_ & new_G1926_ & new_G3795_;
  assign new_G3846_ = new_G3823_ & new_G1921_ & new_G3795_;
  assign new_G3849_ = new_G3841_ | new_G3839_ | new_G3840_;
  assign new_G3960_ = ~new_G5409_ | ~new_G5412_;
  assign new_G5413_ = ~new_G5409_;
  assign new_G3963_ = ~new_G5417_ | ~new_G5420_;
  assign new_G4010_ = new_G3998_ & new_G1238_ & new_G3972_;
  assign new_G4068_ = new_G4056_ & new_G1916_ & new_G4030_;
  assign new_G4358_ = ~new_G4356_ | ~new_G4357_;
  assign new_G4416_ = ~new_G4414_ | ~new_G4415_;
  assign new_G4480_ = ~new_G4474_;
  assign new_G4483_ = ~new_G4474_ | ~new_G4481_;
  assign new_G4568_ = ~new_G4562_;
  assign new_G4571_ = ~new_G4562_ | ~new_G4569_;
  assign new_G4822_ = ~new_G4820_ | ~new_G4821_;
  assign new_G4880_ = ~new_G4878_ | ~new_G4879_;
  assign new_G4938_ = ~new_G4936_ | ~new_G4937_;
  assign new_G5022_ = ~new_G5016_;
  assign new_G5025_ = ~new_G5016_ | ~new_G5023_;
  assign new_G1258_ = new_G1256_ | new_G1257_;
  assign new_G1263_ = new_G1261_ | new_G1262_;
  assign new_G1268_ = new_G1266_ | new_G1267_;
  assign new_G1273_ = new_G1271_ | new_G1272_;
  assign new_G1936_ = new_G1934_ | new_G1935_;
  assign new_G1944_ = new_G1942_ | new_G1943_;
  assign new_G1949_ = new_G1947_ | new_G1948_;
  assign new_G1954_ = new_G1952_ | new_G1953_;
  assign new_G3536_ = ~new_G5247_ | ~new_G5250_;
  assign new_G3541_ = ~new_G5255_ | ~new_G5258_;
  assign new_G3791_ = new_G3783_ | new_G3781_ | new_G3782_;
  assign new_G3792_ = new_G3786_ | new_G3784_ | new_G3785_;
  assign new_G3793_ = new_G3789_ | new_G3787_ | new_G3788_;
  assign new_G3850_ = new_G3844_ | new_G3842_ | new_G3843_;
  assign new_G3851_ = new_G3847_ | new_G3845_ | new_G3846_;
  assign new_G3961_ = ~new_G5406_ | ~new_G5413_;
  assign new_G3965_ = ~new_G3963_ | ~new_G3964_;
  assign new_G4024_ = new_G4011_ | new_G4009_ | new_G4010_;
  assign new_G4082_ = new_G4069_ | new_G4067_ | new_G4068_;
  assign new_G4482_ = ~new_G4477_ | ~new_G4480_;
  assign new_G4570_ = ~new_G4565_ | ~new_G4568_;
  assign new_G5024_ = ~new_G5019_ | ~new_G5022_;
  assign new_G1666_ = new_G1645_ & new_G3790_ & new_G1609_;
  assign new_G1670_ = new_G1645_ & new_G3849_ & new_G1621_;
  assign new_G2337_ = new_G2316_ & new_G3790_ & new_G2281_;
  assign new_G2341_ = new_G2316_ & new_G3849_ & new_G2293_;
  assign new_G719_ = new_G2454_ & new_G3790_ & new_G2418_;
  assign new_G758_ = new_G2454_ & new_G3849_ & new_G2430_;
  assign new_G798_ = new_G2512_ & new_G3849_ & new_G2488_;
  assign G838 = ~new_G3849_;
  assign new_G856_ = new_G2512_ & new_G3790_ & new_G2476_;
  assign G861 = ~new_G3790_;
  assign new_G3538_ = ~new_G3536_ | ~new_G3537_;
  assign new_G3543_ = ~new_G3541_ | ~new_G3542_;
  assign new_G3962_ = ~new_G3960_ | ~new_G3961_;
  assign new_G4364_ = ~new_G4358_;
  assign new_G4367_ = ~new_G4358_ | ~new_G4365_;
  assign new_G4422_ = ~new_G4416_;
  assign new_G4425_ = ~new_G4416_ | ~new_G4423_;
  assign new_G4484_ = ~new_G4482_ | ~new_G4483_;
  assign new_G4572_ = ~new_G4570_ | ~new_G4571_;
  assign new_G4828_ = ~new_G4822_;
  assign new_G4831_ = ~new_G4822_ | ~new_G4829_;
  assign new_G4886_ = ~new_G4880_;
  assign new_G4889_ = ~new_G4880_ | ~new_G4887_;
  assign new_G4944_ = ~new_G4938_;
  assign new_G4947_ = ~new_G4938_ | ~new_G4945_;
  assign new_G5026_ = ~new_G5024_ | ~new_G5025_;
  assign new_G571_ = ~new_G1273_;
  assign new_G572_ = ~new_G1268_;
  assign new_G573_ = ~new_G1263_;
  assign new_G574_ = ~new_G1258_;
  assign new_G581_ = ~new_G1954_;
  assign new_G582_ = ~new_G1949_;
  assign new_G583_ = ~new_G1944_;
  assign new_G584_ = ~new_G1936_;
  assign G623 = ~new_G1936_;
  assign new_G1576_ = new_G1564_ & new_G4082_ & new_G1540_;
  assign new_G1578_ = new_G1564_ & new_G4024_ & new_G1528_;
  assign new_G659_ = new_G1668_ | new_G1667_ | new_G1664_ | new_G1666_;
  assign new_G1672_ = new_G1645_ & new_G3791_ & new_G1609_;
  assign new_G1676_ = new_G1645_ & new_G3850_ & new_G1621_;
  assign new_G1678_ = new_G1645_ & new_G3792_ & new_G1609_;
  assign new_G1682_ = new_G1645_ & new_G3851_ & new_G1621_;
  assign new_G1684_ = new_G1645_ & new_G3793_ & new_G1609_;
  assign new_G2250_ = new_G2238_ & new_G4082_ & new_G2215_;
  assign new_G2252_ = new_G2238_ & new_G4024_ & new_G2203_;
  assign new_G691_ = new_G2339_ | new_G2338_ | new_G2335_ | new_G2337_;
  assign new_G2343_ = new_G2316_ & new_G3791_ & new_G2281_;
  assign new_G2347_ = new_G2316_ & new_G3850_ & new_G2293_;
  assign new_G2349_ = new_G2316_ & new_G3792_ & new_G2281_;
  assign new_G2353_ = new_G2316_ & new_G3851_ & new_G2293_;
  assign new_G2355_ = new_G2316_ & new_G3793_ & new_G2281_;
  assign G722 = new_G721_ | new_G720_ | new_G718_ | new_G719_;
  assign new_G743_ = new_G3594_ & new_G4082_ & new_G3570_;
  assign new_G744_ = new_G3594_ & new_G4024_ & new_G3558_;
  assign new_G748_ = new_G2454_ & new_G3851_ & new_G2430_;
  assign new_G749_ = new_G2454_ & new_G3793_ & new_G2418_;
  assign new_G753_ = new_G2454_ & new_G3850_ & new_G2430_;
  assign new_G754_ = new_G2454_ & new_G3792_ & new_G2418_;
  assign new_G759_ = new_G2454_ & new_G3791_ & new_G2418_;
  assign new_G783_ = new_G3696_ & new_G4082_ & new_G3672_;
  assign new_G784_ = new_G3696_ & new_G4024_ & new_G3660_;
  assign new_G788_ = new_G2512_ & new_G3851_ & new_G2488_;
  assign new_G789_ = new_G2512_ & new_G3793_ & new_G2476_;
  assign new_G793_ = new_G2512_ & new_G3850_ & new_G2488_;
  assign new_G794_ = new_G2512_ & new_G3792_ & new_G2476_;
  assign new_G799_ = new_G2512_ & new_G3791_ & new_G2476_;
  assign new_G3735_ = G3717 & new_G1936_ & G3724;
  assign G832 = ~new_G4082_;
  assign G834 = ~new_G3851_;
  assign G836 = ~new_G3850_;
  assign new_G3835_ = ~new_G3965_;
  assign G859 = new_G858_ | new_G857_ | new_G855_ | new_G856_;
  assign G871 = ~new_G4024_;
  assign G873 = ~new_G3793_;
  assign G875 = ~new_G3792_;
  assign G877 = ~new_G3791_;
  assign G998 = new_G3538_;
  assign G1000 = new_G3543_;
  assign new_G3651_ = new_G3965_ & new_G3632_;
  assign new_G4013_ = new_G3998_ & new_G1273_ & new_G3972_;
  assign new_G4016_ = new_G3998_ & new_G1268_ & new_G3972_;
  assign new_G4019_ = new_G3998_ & new_G1263_ & new_G3972_;
  assign new_G4022_ = new_G3998_ & new_G1258_ & new_G3972_;
  assign new_G4071_ = new_G4056_ & new_G1954_ & new_G4030_;
  assign new_G4074_ = new_G4056_ & new_G1949_ & new_G4030_;
  assign new_G4077_ = new_G4056_ & new_G1944_ & new_G4030_;
  assign new_G4080_ = new_G4056_ & new_G1936_ & new_G4030_;
  assign new_G4096_ = ~new_G4113_ | ~new_G1936_;
  assign new_G4366_ = ~new_G4361_ | ~new_G4364_;
  assign new_G4424_ = ~new_G4419_ | ~new_G4422_;
  assign new_G4830_ = ~new_G4825_ | ~new_G4828_;
  assign new_G4888_ = ~new_G4883_ | ~new_G4886_;
  assign new_G4946_ = ~new_G4941_ | ~new_G4944_;
  assign G575 = new_G574_ & new_G573_ & new_G572_ & new_G571_ & new_G570_ & new_G569_ & new_G568_ & new_G566_ & new_G567_;
  assign G585 = new_G584_ & new_G583_ & new_G582_ & new_G581_ & new_G580_ & new_G579_ & new_G578_ & new_G576_ & new_G577_;
  assign new_G640_ = new_G1580_ | new_G1579_ | new_G1576_ | new_G1578_;
  assign G661 = new_G659_ & new_G1606_;
  assign new_G662_ = new_G1674_ | new_G1673_ | new_G1670_ | new_G1672_;
  assign new_G665_ = new_G1680_ | new_G1679_ | new_G1676_ | new_G1678_;
  assign new_G668_ = new_G1686_ | new_G1685_ | new_G1682_ | new_G1684_;
  assign new_G674_ = new_G2254_ | new_G2253_ | new_G2250_ | new_G2252_;
  assign G693 = new_G691_ & new_G2279_;
  assign new_G694_ = new_G2345_ | new_G2344_ | new_G2341_ | new_G2343_;
  assign new_G697_ = new_G2351_ | new_G2350_ | new_G2347_ | new_G2349_;
  assign new_G700_ = new_G2357_ | new_G2356_ | new_G2353_ | new_G2355_;
  assign G747 = new_G746_ | new_G745_ | new_G743_ | new_G744_;
  assign G752 = new_G751_ | new_G750_ | new_G748_ | new_G749_;
  assign G757 = new_G756_ | new_G755_ | new_G753_ | new_G754_;
  assign G762 = new_G761_ | new_G760_ | new_G758_ | new_G759_;
  assign G787 = new_G786_ | new_G785_ | new_G783_ | new_G784_;
  assign G792 = new_G791_ | new_G790_ | new_G788_ | new_G789_;
  assign G797 = new_G796_ | new_G795_ | new_G793_ | new_G794_;
  assign G802 = new_G801_ | new_G800_ | new_G798_ | new_G799_;
  assign new_G817_ = new_G3735_ | new_G3734_ | new_G3731_ | new_G3733_;
  assign new_G839_ = new_G3823_ & new_G3835_ & new_G3803_;
  assign new_G3540_ = ~new_G3538_;
  assign new_G3545_ = ~new_G3543_;
  assign new_G3777_ = ~new_G3962_;
  assign new_G3648_ = new_G3962_ & new_G3632_;
  assign new_G4025_ = new_G4014_ | new_G4012_ | new_G4013_;
  assign new_G4026_ = new_G4017_ | new_G4015_ | new_G4016_;
  assign new_G4027_ = new_G4020_ | new_G4018_ | new_G4019_;
  assign new_G4028_ = new_G4023_ | new_G4021_ | new_G4022_;
  assign new_G4083_ = new_G4072_ | new_G4070_ | new_G4071_;
  assign new_G4084_ = new_G4075_ | new_G4073_ | new_G4074_;
  assign new_G4085_ = new_G4078_ | new_G4076_ | new_G4077_;
  assign new_G4086_ = new_G4081_ | new_G4079_ | new_G4080_;
  assign new_G4368_ = ~new_G4366_ | ~new_G4367_;
  assign new_G4426_ = ~new_G4424_ | ~new_G4425_;
  assign new_G4490_ = ~new_G4484_;
  assign new_G4493_ = ~new_G4484_ | ~new_G4491_;
  assign new_G4578_ = ~new_G4572_;
  assign new_G4581_ = ~new_G4572_ | ~new_G4579_;
  assign new_G4832_ = ~new_G4830_ | ~new_G4831_;
  assign new_G4890_ = ~new_G4888_ | ~new_G4889_;
  assign new_G4948_ = ~new_G4946_ | ~new_G4947_;
  assign new_G5032_ = ~new_G5026_;
  assign new_G5035_ = ~new_G5026_ | ~new_G5033_;
  assign G642 = new_G640_ & new_G1526_;
  assign G664 = new_G662_ & new_G1606_;
  assign G667 = new_G665_ & new_G1606_;
  assign G670 = new_G668_ & new_G1606_;
  assign G676 = new_G674_ & new_G2202_;
  assign G696 = new_G694_ & new_G2279_;
  assign G699 = new_G697_ & new_G2279_;
  assign G702 = new_G700_ & new_G2279_;
  assign new_G811_ = new_G4113_ & new_G4096_;
  assign new_G812_ = new_G4096_ & new_G1936_;
  assign G818 = new_G816_ & new_G817_;
  assign new_G853_ = new_G3970_ & new_G3535_ & new_G3545_ & G562 & new_G3540_;
  assign new_G878_ = new_G3765_ & new_G3777_ & new_G3745_;
  assign new_G4492_ = ~new_G4487_ | ~new_G4490_;
  assign new_G4580_ = ~new_G4575_ | ~new_G4578_;
  assign new_G5034_ = ~new_G5029_ | ~new_G5032_;
  assign new_G1582_ = new_G1564_ & new_G4083_ & new_G1540_;
  assign new_G1584_ = new_G1564_ & new_G4025_ & new_G1528_;
  assign new_G1588_ = new_G1564_ & new_G4084_ & new_G1540_;
  assign new_G1590_ = new_G1564_ & new_G4026_ & new_G1528_;
  assign new_G1594_ = new_G1564_ & new_G4085_ & new_G1540_;
  assign new_G1596_ = new_G1564_ & new_G4027_ & new_G1528_;
  assign new_G1600_ = new_G1564_ & new_G4086_ & new_G1540_;
  assign new_G1602_ = new_G1564_ & new_G4028_ & new_G1528_;
  assign new_G2256_ = new_G2238_ & new_G4083_ & new_G2215_;
  assign new_G2258_ = new_G2238_ & new_G4025_ & new_G2203_;
  assign new_G2262_ = new_G2238_ & new_G4084_ & new_G2215_;
  assign new_G2264_ = new_G2238_ & new_G4026_ & new_G2203_;
  assign new_G2268_ = new_G2238_ & new_G4085_ & new_G2215_;
  assign new_G2270_ = new_G2238_ & new_G4027_ & new_G2203_;
  assign new_G2274_ = new_G2238_ & new_G4086_ & new_G2215_;
  assign new_G2276_ = new_G2238_ & new_G4028_ & new_G2203_;
  assign new_G708_ = new_G3696_ & new_G4086_ & new_G3672_;
  assign new_G709_ = new_G3696_ & new_G4028_ & new_G3660_;
  assign new_G723_ = new_G3594_ & new_G4086_ & new_G3570_;
  assign new_G724_ = new_G3594_ & new_G4028_ & new_G3558_;
  assign new_G728_ = new_G3594_ & new_G4085_ & new_G3570_;
  assign new_G729_ = new_G3594_ & new_G4027_ & new_G3558_;
  assign new_G733_ = new_G3594_ & new_G4084_ & new_G3570_;
  assign new_G734_ = new_G3594_ & new_G4026_ & new_G3558_;
  assign new_G738_ = new_G3594_ & new_G4083_ & new_G3570_;
  assign new_G739_ = new_G3594_ & new_G4025_ & new_G3558_;
  assign new_G768_ = new_G3696_ & new_G4085_ & new_G3672_;
  assign new_G769_ = new_G3696_ & new_G4027_ & new_G3660_;
  assign new_G773_ = new_G3696_ & new_G4084_ & new_G3672_;
  assign new_G774_ = new_G3696_ & new_G4026_ & new_G3660_;
  assign new_G778_ = new_G3696_ & new_G4083_ & new_G3672_;
  assign new_G779_ = new_G3696_ & new_G4025_ & new_G3660_;
  assign G813 = new_G811_ | new_G812_;
  assign G824 = ~new_G4086_;
  assign G826 = ~new_G4085_;
  assign G828 = ~new_G4084_;
  assign G830 = ~new_G4083_;
  assign G854 = G245 & new_G852_ & new_G853_;
  assign G863 = ~new_G4028_;
  assign G865 = ~new_G4027_;
  assign G867 = ~new_G4026_;
  assign G869 = ~new_G4025_;
  assign new_G4374_ = ~new_G4368_;
  assign new_G4377_ = ~new_G4368_ | ~new_G4375_;
  assign new_G4432_ = ~new_G4426_;
  assign new_G4435_ = ~new_G4426_ | ~new_G4433_;
  assign new_G4494_ = ~new_G4492_ | ~new_G4493_;
  assign new_G4582_ = ~new_G4580_ | ~new_G4581_;
  assign new_G4838_ = ~new_G4832_;
  assign new_G4841_ = ~new_G4832_ | ~new_G4839_;
  assign new_G4896_ = ~new_G4890_;
  assign new_G4899_ = ~new_G4890_ | ~new_G4897_;
  assign new_G4954_ = ~new_G4948_;
  assign new_G4957_ = ~new_G4948_ | ~new_G4955_;
  assign new_G5036_ = ~new_G5034_ | ~new_G5035_;
  assign new_G643_ = new_G1586_ | new_G1585_ | new_G1582_ | new_G1584_;
  assign new_G646_ = new_G1592_ | new_G1591_ | new_G1588_ | new_G1590_;
  assign new_G649_ = new_G1598_ | new_G1597_ | new_G1594_ | new_G1596_;
  assign new_G652_ = new_G1604_ | new_G1603_ | new_G1600_ | new_G1602_;
  assign new_G677_ = new_G2260_ | new_G2259_ | new_G2256_ | new_G2258_;
  assign new_G680_ = new_G2266_ | new_G2265_ | new_G2262_ | new_G2264_;
  assign new_G683_ = new_G2272_ | new_G2271_ | new_G2268_ | new_G2270_;
  assign new_G686_ = new_G2278_ | new_G2277_ | new_G2274_ | new_G2276_;
  assign G712 = new_G711_ | new_G710_ | new_G708_ | new_G709_;
  assign G727 = new_G726_ | new_G725_ | new_G723_ | new_G724_;
  assign G732 = new_G731_ | new_G730_ | new_G728_ | new_G729_;
  assign G737 = new_G736_ | new_G735_ | new_G733_ | new_G734_;
  assign G742 = new_G741_ | new_G740_ | new_G738_ | new_G739_;
  assign G772 = new_G771_ | new_G770_ | new_G768_ | new_G769_;
  assign G777 = new_G776_ | new_G775_ | new_G773_ | new_G774_;
  assign G782 = new_G781_ | new_G780_ | new_G778_ | new_G779_;
  assign new_G4376_ = ~new_G4371_ | ~new_G4374_;
  assign new_G4434_ = ~new_G4429_ | ~new_G4432_;
  assign new_G4840_ = ~new_G4835_ | ~new_G4838_;
  assign new_G4898_ = ~new_G4893_ | ~new_G4896_;
  assign new_G4956_ = ~new_G4951_ | ~new_G4954_;
  assign G645 = new_G643_ & new_G1526_;
  assign G648 = new_G646_ & new_G1526_;
  assign G651 = new_G649_ & new_G1526_;
  assign G654 = new_G652_ & new_G1526_;
  assign G679 = new_G677_ & new_G2202_;
  assign G682 = new_G680_ & new_G2202_;
  assign G685 = new_G683_ & new_G2202_;
  assign G688 = new_G686_ & new_G2202_;
  assign new_G4378_ = ~new_G4376_ | ~new_G4377_;
  assign new_G4436_ = ~new_G4434_ | ~new_G4435_;
  assign new_G4500_ = ~new_G4494_;
  assign new_G4503_ = ~new_G4494_ | ~new_G4501_;
  assign new_G4588_ = ~new_G4582_;
  assign new_G4591_ = ~new_G4582_ | ~new_G4589_;
  assign new_G4842_ = ~new_G4840_ | ~new_G4841_;
  assign new_G4900_ = ~new_G4898_ | ~new_G4899_;
  assign new_G4958_ = ~new_G4956_ | ~new_G4957_;
  assign new_G5042_ = ~new_G5036_;
  assign new_G5045_ = ~new_G5036_ | ~new_G5043_;
  assign new_G4502_ = ~new_G4497_ | ~new_G4500_;
  assign new_G4590_ = ~new_G4585_ | ~new_G4588_;
  assign new_G5044_ = ~new_G5039_ | ~new_G5042_;
  assign new_G4384_ = ~new_G4378_;
  assign new_G4387_ = ~new_G4378_ | ~new_G4385_;
  assign new_G4442_ = ~new_G4436_;
  assign new_G4445_ = ~new_G4436_ | ~new_G4443_;
  assign new_G4504_ = ~new_G4502_ | ~new_G4503_;
  assign new_G4592_ = ~new_G4590_ | ~new_G4591_;
  assign new_G4848_ = ~new_G4842_;
  assign new_G4851_ = ~new_G4842_ | ~new_G4849_;
  assign new_G4906_ = ~new_G4900_;
  assign new_G4909_ = ~new_G4900_ | ~new_G4907_;
  assign new_G4964_ = ~new_G4958_;
  assign new_G4967_ = ~new_G4958_ | ~new_G4965_;
  assign new_G5046_ = ~new_G5044_ | ~new_G5045_;
  assign new_G4386_ = ~new_G4381_ | ~new_G4384_;
  assign new_G4444_ = ~new_G4439_ | ~new_G4442_;
  assign new_G4850_ = ~new_G4845_ | ~new_G4848_;
  assign new_G4908_ = ~new_G4903_ | ~new_G4906_;
  assign new_G4966_ = ~new_G4961_ | ~new_G4964_;
  assign new_G4388_ = ~new_G4386_ | ~new_G4387_;
  assign new_G4446_ = ~new_G4444_ | ~new_G4445_;
  assign new_G4510_ = ~new_G4504_;
  assign new_G4513_ = ~new_G4504_ | ~new_G4511_;
  assign new_G4598_ = ~new_G4592_;
  assign new_G4601_ = ~new_G4592_ | ~new_G4599_;
  assign new_G4852_ = ~new_G4850_ | ~new_G4851_;
  assign new_G4910_ = ~new_G4908_ | ~new_G4909_;
  assign new_G4968_ = ~new_G4966_ | ~new_G4967_;
  assign new_G5052_ = ~new_G5046_;
  assign new_G5055_ = ~new_G5046_ | ~new_G5053_;
  assign new_G4512_ = ~new_G4507_ | ~new_G4510_;
  assign new_G4600_ = ~new_G4595_ | ~new_G4598_;
  assign new_G5054_ = ~new_G5049_ | ~new_G5052_;
  assign new_G4394_ = ~new_G4388_;
  assign new_G4397_ = ~new_G4388_ | ~new_G4395_;
  assign new_G4452_ = ~new_G4446_;
  assign new_G4455_ = ~new_G4446_ | ~new_G4453_;
  assign new_G4514_ = ~new_G4512_ | ~new_G4513_;
  assign new_G4602_ = ~new_G4600_ | ~new_G4601_;
  assign new_G4858_ = ~new_G4852_;
  assign new_G4861_ = ~new_G4852_ | ~new_G4859_;
  assign new_G4916_ = ~new_G4910_;
  assign new_G4919_ = ~new_G4910_ | ~new_G4917_;
  assign new_G4974_ = ~new_G4968_;
  assign new_G4977_ = ~new_G4968_ | ~new_G4975_;
  assign new_G5056_ = ~new_G5054_ | ~new_G5055_;
  assign new_G4396_ = ~new_G4391_ | ~new_G4394_;
  assign new_G4454_ = ~new_G4449_ | ~new_G4452_;
  assign new_G4860_ = ~new_G4855_ | ~new_G4858_;
  assign new_G4918_ = ~new_G4913_ | ~new_G4916_;
  assign new_G4976_ = ~new_G4971_ | ~new_G4974_;
  assign new_G4398_ = ~new_G4396_ | ~new_G4397_;
  assign new_G4456_ = ~new_G4454_ | ~new_G4455_;
  assign new_G4520_ = ~new_G4514_;
  assign new_G4523_ = ~new_G4514_ | ~new_G4521_;
  assign new_G4608_ = ~new_G4602_;
  assign new_G4611_ = ~new_G4602_ | ~new_G4609_;
  assign new_G4862_ = ~new_G4860_ | ~new_G4861_;
  assign new_G4920_ = ~new_G4918_ | ~new_G4919_;
  assign new_G4978_ = ~new_G4976_ | ~new_G4977_;
  assign new_G5062_ = ~new_G5056_;
  assign new_G5065_ = ~new_G5056_ | ~new_G5063_;
  assign new_G4522_ = ~new_G4517_ | ~new_G4520_;
  assign new_G4610_ = ~new_G4605_ | ~new_G4608_;
  assign new_G5064_ = ~new_G5059_ | ~new_G5062_;
  assign new_G4404_ = ~new_G4398_;
  assign new_G1488_ = ~new_G4398_ | ~new_G4405_;
  assign new_G4462_ = ~new_G4456_;
  assign new_G1493_ = ~new_G4456_ | ~new_G4463_;
  assign new_G4868_ = ~new_G4862_;
  assign new_G2165_ = ~new_G4862_ | ~new_G4869_;
  assign new_G4926_ = ~new_G4920_;
  assign new_G2170_ = ~new_G4920_ | ~new_G4927_;
  assign new_G4524_ = ~new_G4522_ | ~new_G4523_;
  assign new_G4612_ = ~new_G4610_ | ~new_G4611_;
  assign new_G4984_ = ~new_G4978_;
  assign new_G4987_ = ~new_G4978_ | ~new_G4985_;
  assign new_G5066_ = ~new_G5064_ | ~new_G5065_;
  assign new_G1487_ = ~new_G4401_ | ~new_G4404_;
  assign new_G1492_ = ~new_G4459_ | ~new_G4462_;
  assign new_G2164_ = ~new_G4865_ | ~new_G4868_;
  assign new_G2169_ = ~new_G4923_ | ~new_G4926_;
  assign new_G4986_ = ~new_G4981_ | ~new_G4984_;
  assign new_G1489_ = ~new_G1487_ | ~new_G1488_;
  assign new_G1494_ = ~new_G1492_ | ~new_G1493_;
  assign new_G2166_ = ~new_G2164_ | ~new_G2165_;
  assign new_G2171_ = ~new_G2169_ | ~new_G2170_;
  assign new_G4530_ = ~new_G4524_;
  assign new_G4533_ = ~new_G4524_ | ~new_G4531_;
  assign new_G4618_ = ~new_G4612_;
  assign new_G4543_ = ~new_G4612_ | ~new_G4619_;
  assign new_G4988_ = ~new_G4986_ | ~new_G4987_;
  assign new_G5072_ = ~new_G5066_;
  assign new_G4997_ = ~new_G5066_ | ~new_G5073_;
  assign new_G4532_ = ~new_G4527_ | ~new_G4530_;
  assign new_G4542_ = ~new_G4615_ | ~new_G4618_;
  assign new_G4996_ = ~new_G5069_ | ~new_G5072_;
  assign new_G1513_ = new_G1502_ & new_G1494_ & new_G1462_;
  assign new_G1514_ = new_G1502_ & new_G1489_ & new_G1458_;
  assign new_G1515_ = G1497 & new_G1494_ & new_G1483_;
  assign new_G1516_ = G1497 & new_G1489_ & new_G1486_;
  assign new_G4994_ = ~new_G4988_;
  assign new_G2184_ = ~new_G4988_ | ~new_G4995_;
  assign new_G2190_ = new_G2179_ & new_G2171_ & new_G2139_;
  assign new_G2191_ = new_G2179_ & new_G2166_ & new_G2135_;
  assign new_G2192_ = G2174 & new_G2171_ & new_G2160_;
  assign new_G2193_ = G2174 & new_G2166_ & new_G2163_;
  assign new_G4534_ = ~new_G4532_ | ~new_G4533_;
  assign new_G4544_ = ~new_G4542_ | ~new_G4543_;
  assign new_G4998_ = ~new_G4996_ | ~new_G4997_;
  assign new_G2183_ = ~new_G4991_ | ~new_G4994_;
  assign new_G4620_ = new_G1516_ | new_G1515_ | new_G1513_ | new_G1514_;
  assign new_G5074_ = new_G2193_ | new_G2192_ | new_G2190_ | new_G2191_;
  assign new_G4540_ = ~new_G4534_;
  assign new_G1507_ = ~new_G4534_ | ~new_G4541_;
  assign new_G4550_ = ~new_G4544_;
  assign new_G1510_ = ~new_G4544_ | ~new_G4551_;
  assign new_G2185_ = ~new_G2183_ | ~new_G2184_;
  assign new_G5004_ = ~new_G4998_;
  assign new_G2187_ = ~new_G4998_ | ~new_G5005_;
  assign new_G1506_ = ~new_G4537_ | ~new_G4540_;
  assign new_G1509_ = ~new_G4547_ | ~new_G4550_;
  assign new_G4626_ = ~new_G4620_;
  assign new_G2186_ = ~new_G5001_ | ~new_G5004_;
  assign new_G2195_ = G2174 & new_G2185_;
  assign new_G5080_ = ~new_G5074_;
  assign new_G1508_ = ~new_G1506_ | ~new_G1507_;
  assign new_G1511_ = ~new_G1509_ | ~new_G1510_;
  assign new_G2188_ = ~new_G2186_ | ~new_G2187_;
  assign new_G1512_ = ~new_G1511_;
  assign new_G1518_ = G1497 & new_G1508_;
  assign new_G2189_ = ~new_G2188_;
  assign new_G1517_ = new_G1512_ & new_G1502_;
  assign new_G2194_ = new_G2189_ & new_G2179_;
  assign new_G4623_ = new_G1517_ | new_G1518_;
  assign new_G5077_ = new_G2194_ | new_G2195_;
  assign new_G1519_ = ~new_G4623_ | ~new_G4626_;
  assign new_G4627_ = ~new_G4623_;
  assign new_G2196_ = ~new_G5077_ | ~new_G5080_;
  assign new_G5081_ = ~new_G5077_;
  assign new_G1520_ = ~new_G4620_ | ~new_G4627_;
  assign new_G2197_ = ~new_G5074_ | ~new_G5081_;
  assign new_G1521_ = ~new_G1519_ | ~new_G1520_;
  assign new_G2198_ = ~new_G2196_ | ~new_G2197_;
  assign new_G840_ = new_G3823_ & new_G2198_ & new_G3795_;
  assign new_G879_ = new_G3765_ & new_G1521_ & new_G3737_;
  assign new_G1524_ = ~new_G1521_;
  assign new_G2201_ = ~new_G2198_;
  assign G843 = new_G842_ | new_G841_ | new_G839_ | new_G840_;
  assign G882 = new_G881_ | new_G880_ | new_G878_ | new_G879_;
  assign new_G3649_ = new_G1524_ & new_G3628_;
  assign new_G3652_ = new_G2201_ & new_G3628_;
  assign new_G3657_ = new_G3648_ | new_G3649_;
  assign new_G3658_ = new_G3651_ | new_G3652_;
  assign new_G3636_ = new_G3657_ & new_G3622_;
  assign new_G3639_ = new_G3658_ & new_G3622_;
  assign new_G3642_ = new_G3657_ & new_G3622_;
  assign new_G3645_ = new_G3658_ & new_G3622_;
  assign new_G3653_ = new_G3636_ | new_G3637_;
  assign new_G3654_ = new_G3639_ | new_G3640_;
  assign new_G3655_ = new_G3642_ | new_G3643_;
  assign new_G3656_ = new_G3645_ | new_G3646_;
  assign new_G763_ = new_G2454_ & new_G3656_ & new_G2430_;
  assign new_G764_ = new_G2454_ & new_G3655_ & new_G2418_;
  assign new_G803_ = new_G2512_ & new_G3656_ & new_G2488_;
  assign new_G804_ = new_G2512_ & new_G3655_ & new_G2476_;
  assign new_G1657_ = new_G1645_ & new_G3654_ & new_G1621_;
  assign new_G1659_ = new_G1645_ & new_G3653_ & new_G1609_;
  assign new_G2328_ = new_G2316_ & new_G3654_ & new_G2293_;
  assign new_G2330_ = new_G2316_ & new_G3653_ & new_G2281_;
  assign new_G1662_ = new_G1661_ | new_G1660_ | new_G1657_ | new_G1659_;
  assign new_G2333_ = new_G2332_ | new_G2331_ | new_G2328_ | new_G2330_;
  assign G767 = new_G766_ | new_G765_ | new_G763_ | new_G764_;
  assign G807 = new_G806_ | new_G805_ | new_G803_ | new_G804_;
  assign new_G657_ = new_G1662_ & new_G1606_;
  assign new_G689_ = new_G2333_ & new_G2279_;
  assign G658 = ~new_G657_;
  assign G690 = ~new_G689_;
endmodule


