// NOR_NOT mapped module c1355

module c1355 (
  input  G1gat   ,
  input  G8gat   ,
  input  G15gat  ,
  input  G22gat  ,
  input  G29gat  ,
  input  G36gat  ,
  input  G43gat  ,
  input  G50gat  ,
  input  G57gat  ,
  input  G64gat  ,
  input  G71gat  ,
  input  G78gat  ,
  input  G85gat  ,
  input  G92gat  ,
  input  G99gat  ,
  input  G106gat ,
  input  G113gat ,
  input  G120gat ,
  input  G127gat ,
  input  G134gat ,
  input  G141gat ,
  input  G148gat ,
  input  G155gat ,
  input  G162gat ,
  input  G169gat ,
  input  G176gat ,
  input  G183gat ,
  input  G190gat ,
  input  G197gat ,
  input  G204gat ,
  input  G211gat ,
  input  G218gat ,
  input  G225gat ,
  input  G226gat ,
  input  G227gat ,
  input  G228gat ,
  input  G229gat ,
  input  G230gat ,
  input  G231gat ,
  input  G232gat ,
  input  G233gat ,
  output G1324gat,
  output G1325gat,
  output G1326gat,
  output G1327gat,
  output G1328gat,
  output G1329gat,
  output G1330gat,
  output G1331gat,
  output G1332gat,
  output G1333gat,
  output G1334gat,
  output G1335gat,
  output G1336gat,
  output G1337gat,
  output G1338gat,
  output G1339gat,
  output G1340gat,
  output G1341gat,
  output G1342gat,
  output G1343gat,
  output G1344gat,
  output G1345gat,
  output G1346gat,
  output G1347gat,
  output G1348gat,
  output G1349gat,
  output G1350gat,
  output G1351gat,
  output G1352gat,
  output G1353gat,
  output G1354gat,
  output G1355gat);

  wire wr_33;
  wire wr_34;
  wire wr_35;
  wire wr_36;
  wire wr_37;
  wire wr_38;
  wire wr_39;
  wire wr_40;
  wire wr_41;
  wire wr_42;
  wire wr_43;
  wire wr_44;
  wire wr_45;
  wire wr_46;
  wire wr_47;
  wire wr_48;
  wire wr_49;
  wire wr_50;
  wire wr_51;
  wire wr_52;
  wire wr_53;
  wire wr_54;
  wire wr_55;
  wire wr_56;
  wire wr_57;
  wire wr_58;
  wire wr_59;
  wire wr_60;
  wire wr_61;
  wire wr_62;
  wire wr_63;
  wire wr_64;
  wire wr_65;
  wire wr_66;
  wire wr_67;
  wire wr_68;
  wire wr_69;
  wire wr_70;
  wire wr_71;
  wire wr_72;
  wire wr_73;
  wire wr_74;
  wire wr_75;
  wire wr_76;
  wire wr_77;
  wire wr_78;
  wire wr_79;
  wire wr_80;
  wire wr_81;
  wire wr_82;
  wire wr_83;
  wire wr_84;
  wire wr_85;
  wire wr_86;
  wire wr_87;
  wire wr_88;
  wire wr_89;
  wire wr_90;
  wire wr_91;
  wire wr_92;
  wire wr_93;
  wire wr_94;
  wire wr_95;
  wire wr_96;
  wire wr_97;
  wire wr_98;
  wire wr_99;
  wire wr_100;
  wire wr_101;
  wire wr_102;
  wire wr_103;
  wire wr_104;
  wire wr_105;
  wire wr_106;
  wire wr_107;
  wire wr_108;
  wire wr_109;
  wire wr_110;
  wire wr_111;
  wire wr_112;
  wire wr_113;
  wire wr_114;
  wire wr_115;
  wire wr_116;
  wire wr_117;
  wire wr_118;
  wire wr_119;
  wire wr_120;
  wire wr_121;
  wire wr_122;
  wire wr_123;
  wire wr_124;
  wire wr_125;
  wire wr_126;
  wire wr_127;
  wire wr_128;
  wire wr_129;
  wire wr_130;
  wire wr_131;
  wire wr_132;
  wire wr_133;
  wire wr_134;
  wire wr_135;
  wire wr_136;
  wire wr_137;
  wire wr_138;
  wire wr_139;
  wire wr_140;
  wire wr_141;
  wire wr_142;
  wire wr_143;
  wire wr_144;
  wire wr_145;
  wire wr_146;
  wire wr_147;
  wire wr_148;
  wire wr_149;
  wire wr_150;
  wire wr_151;
  wire wr_152;
  wire wr_153;
  wire wr_154;
  wire wr_155;
  wire wr_156;
  wire wr_157;
  wire wr_158;
  wire wr_159;
  wire wr_160;
  wire wr_161;
  wire wr_162;
  wire wr_163;
  wire wr_164;
  wire wr_165;
  wire wr_166;
  wire wr_167;
  wire wr_168;
  wire wr_169;
  wire wr_170;
  wire wr_171;
  wire wr_172;
  wire wr_173;
  wire wr_174;
  wire wr_175;
  wire wr_176;
  wire wr_177;
  wire wr_178;
  wire wr_179;
  wire wr_180;
  wire wr_181;
  wire wr_182;
  wire wr_183;
  wire wr_184;
  wire wr_185;
  wire wr_186;
  wire wr_187;
  wire wr_188;
  wire wr_189;
  wire wr_190;
  wire wr_191;
  wire wr_192;
  wire wr_193;
  wire wr_194;
  wire wr_195;
  wire wr_196;
  wire wr_197;
  wire wr_198;
  wire wr_199;
  wire wr_200;
  wire wr_201;
  wire wr_202;
  wire wr_203;
  wire wr_204;
  wire wr_205;
  wire wr_206;
  wire wr_207;
  wire wr_208;
  wire wr_209;
  wire wr_210;
  wire wr_211;
  wire wr_212;
  wire wr_213;
  wire wr_214;
  wire wr_215;
  wire wr_216;
  wire wr_217;
  wire wr_218;
  wire wr_219;
  wire wr_220;
  wire wr_221;
  wire wr_222;
  wire wr_223;
  wire wr_224;
  wire wr_225;
  wire wr_226;
  wire wr_227;
  wire wr_228;
  wire wr_229;
  wire wr_230;
  wire wr_231;
  wire wr_232;
  wire wr_233;
  wire wr_234;
  wire wr_235;
  wire wr_236;
  wire wr_237;
  wire wr_238;
  wire wr_239;
  wire wr_240;
  wire wr_241;
  wire wr_242;
  wire wr_243;
  wire wr_244;
  wire wr_245;
  wire wr_246;
  wire wr_247;
  wire wr_248;
  wire wr_249;
  wire wr_250;
  wire wr_251;
  wire wr_252;
  wire wr_253;
  wire wr_254;
  wire wr_255;
  wire wr_256;
  wire wr_257;
  wire wr_258;
  wire wr_259;
  wire wr_260;
  wire wr_261;
  wire wr_262;
  wire wr_263;
  wire wr_264;
  wire wr_265;
  wire wr_266;
  wire wr_267;
  wire wr_268;
  wire wr_269;
  wire wr_270;
  wire wr_271;
  wire wr_272;
  wire wr_273;
  wire wr_274;
  wire wr_275;
  wire wr_276;
  wire wr_277;
  wire wr_278;
  wire wr_279;
  wire wr_280;
  wire wr_281;
  wire wr_282;
  wire wr_283;
  wire wr_284;
  wire wr_285;
  wire wr_286;
  wire wr_287;
  wire wr_288;
  wire wr_289;
  wire wr_290;
  wire wr_291;
  wire wr_292;
  wire wr_293;
  wire wr_294;
  wire wr_295;
  wire wr_296;
  wire wr_297;
  wire wr_298;
  wire wr_299;
  wire wr_300;
  wire wr_301;
  wire wr_302;
  wire wr_303;
  wire wr_304;
  wire wr_305;
  wire wr_306;
  wire wr_307;
  wire wr_308;
  wire wr_309;
  wire wr_310;
  wire wr_311;
  wire wr_312;
  wire wr_313;
  wire wr_314;
  wire wr_315;
  wire wr_316;
  wire wr_317;
  wire wr_318;
  wire wr_319;
  wire wr_320;
  wire wr_321;
  wire wr_322;
  wire wr_323;
  wire wr_324;
  wire wr_325;
  wire wr_326;
  wire wr_327;
  wire wr_328;
  wire wr_329;
  wire wr_330;
  wire wr_331;
  wire wr_332;
  wire wr_333;
  wire wr_334;
  wire wr_335;
  wire wr_336;
  wire wr_337;
  wire wr_338;
  wire wr_339;
  wire wr_340;
  wire wr_341;
  wire wr_342;
  wire wr_343;
  wire wr_344;
  wire wr_345;
  wire wr_346;
  wire wr_347;
  wire wr_348;
  wire wr_349;
  wire wr_350;
  wire wr_351;
  wire wr_352;
  wire wr_353;
  wire wr_354;
  wire wr_355;
  wire wr_356;
  wire wr_357;
  wire wr_358;
  wire wr_359;
  wire wr_360;
  wire wr_361;
  wire wr_362;
  wire wr_363;
  wire wr_364;
  wire wr_365;
  wire wr_366;
  wire wr_367;
  wire wr_368;
  wire wr_369;
  wire wr_370;
  wire wr_371;
  wire wr_372;
  wire wr_373;
  wire wr_374;
  wire wr_375;
  wire wr_376;
  wire wr_377;
  wire wr_378;
  wire wr_379;
  wire wr_380;
  wire wr_381;
  wire wr_382;
  wire wr_383;
  wire wr_384;
  wire wr_385;
  wire wr_386;
  wire wr_387;
  wire wr_388;
  wire wr_389;
  wire wr_390;
  wire wr_391;
  wire wr_392;
  wire wr_393;
  wire wr_394;
  wire wr_395;
  wire wr_396;
  wire wr_397;
  wire wr_398;
  wire wr_399;
  wire wr_400;
  wire wr_401;
  wire wr_402;
  wire wr_403;
  wire wr_404;
  wire wr_405;
  wire wr_406;
  wire wr_407;
  wire wr_408;
  wire wr_409;
  wire wr_410;
  wire wr_411;
  wire wr_412;
  wire wr_413;
  wire wr_414;
  wire wr_415;
  wire wr_416;
  wire wr_417;
  wire wr_418;
  wire wr_419;
  wire wr_420;
  wire wr_421;
  wire wr_422;
  wire wr_423;
  wire wr_424;
  wire wr_425;
  wire wr_426;
  wire wr_427;
  wire wr_428;
  wire wr_429;
  wire wr_430;
  wire wr_431;
  wire wr_432;
  wire wr_433;
  wire wr_434;
  wire wr_435;
  wire wr_436;
  wire wr_437;
  wire wr_438;
  wire wr_439;
  wire wr_440;
  wire wr_441;
  wire wr_442;
  wire wr_443;
  wire wr_444;
  wire wr_445;
  wire wr_446;
  wire wr_447;
  wire wr_448;
  wire wr_449;
  wire wr_450;
  wire wr_451;
  wire wr_452;
  wire wr_453;
  wire wr_454;
  wire wr_455;
  wire wr_456;
  wire wr_457;
  wire wr_458;
  wire wr_459;
  wire wr_460;
  wire wr_461;
  wire wr_462;
  wire wr_463;
  wire wr_464;
  wire wr_465;
  wire wr_466;
  wire wr_467;
  wire wr_468;
  wire wr_469;
  wire wr_470;
  wire wr_471;
  wire wr_472;
  wire wr_473;
  wire wr_474;
  wire wr_475;
  wire wr_476;
  wire wr_477;
  wire wr_478;
  wire wr_479;
  wire wr_480;
  wire wr_481;
  wire wr_482;
  wire wr_483;
  wire wr_484;
  wire wr_485;
  wire wr_486;
  wire wr_487;
  wire wr_488;
  wire wr_489;
  wire wr_490;
  wire wr_491;
  wire wr_492;
  wire wr_493;
  wire wr_494;
  wire wr_495;
  wire wr_496;
  wire wr_497;
  wire wr_498;
  wire wr_499;
  wire wr_500;
  wire wr_501;
  wire wr_502;
  wire wr_503;
  wire wr_504;
  wire wr_505;
  wire wr_506;
  wire wr_507;
  wire wr_508;
  wire wr_509;
  wire wr_510;
  wire wr_511;
  wire wr_512;
  wire wr_513;
  wire wr_514;
  wire wr_515;
  wire wr_516;
  wire wr_517;
  wire wr_518;
  wire wr_519;
  wire wr_520;
  wire wr_521;
  wire wr_522;
  wire wr_523;
  wire wr_524;
  wire wr_525;
  wire wr_526;
  wire wr_527;
  wire wr_528;
  wire wr_529;
  wire wr_530;
  wire wr_531;
  wire wr_532;
  wire wr_533;
  wire wr_534;
  wire wr_535;
  wire wr_536;
  wire wr_537;
  wire wr_538;
  wire wr_539;
  wire wr_540;
  wire wr_541;
  wire wr_542;
  wire wr_543;
  wire wr_544;
  wire wr_545;
  wire wr_546;
  wire wr_547;
  wire wr_548;
  wire wr_549;
  wire wr_550;
  wire wr_551;
  wire wr_552;
  wire wr_553;
  wire wr_554;
  wire wr_555;
  wire wr_556;
  wire wr_557;
  wire wr_558;
  wire wr_559;
  wire wr_560;
  wire wr_561;
  wire wr_562;
  wire wr_563;
  wire wr_564;
  wire wr_565;
  wire wr_566;
  wire wr_567;
  wire wr_568;
  wire wr_569;
  wire wr_570;
  wire wr_571;
  wire wr_572;
  wire wr_573;
  wire wr_574;
  wire wr_575;
  wire wr_576;
  wire wr_577;
  wire wr_578;
  wire wr_579;
  wire wr_580;
  wire wr_581;
  wire wr_582;
  wire wr_583;
  wire wr_584;
  wire wr_585;
  wire wr_586;
  wire wr_587;
  wire wr_588;
  wire wr_589;
  wire wr_590;
  wire wr_591;
  wire wr_592;
  wire wr_593;
  wire wr_594;
  wire wr_595;
  wire wr_596;
  wire wr_597;
  wire wr_598;
  wire wr_599;
  wire wr_600;
  wire wr_601;
  wire wr_602;
  wire wr_603;
  wire wr_604;
  wire wr_605;
  wire wr_606;
  wire wr_607;
  wire wr_608;
  wire wr_609;
  wire wr_610;
  wire wr_611;
  wire wr_612;
  wire wr_613;
  wire wr_614;
  wire wr_615;
  wire wr_616;
  wire wr_617;
  wire wr_618;
  wire wr_619;
  wire wr_620;
  wire wr_621;
  wire wr_622;
  wire wr_623;
  wire wr_624;
  wire wr_625;
  wire wr_626;
  wire wr_627;
  wire wr_628;
  wire wr_629;
  wire wr_630;
  wire wr_631;

  not    g1( wr_33   ,           G1gat   );
  not    g2( wr_35   ,           G29gat  );
  not    g3( wr_38   ,           G57gat  );
  not    g4( wr_40   ,           G85gat  );
  not    g5( wr_49   ,           G233gat );
  not    g6( wr_52   ,           G113gat );
  not    g7( wr_54   ,           G120gat );
  not    g8( wr_57   ,           G127gat );
  not    g9( wr_59   ,           G134gat );
  not   g10( wr_67   ,           G141gat );
  not   g11( wr_69   ,           G148gat );
  not   g12( wr_72   ,           G155gat );
  not   g13( wr_74   ,           G162gat );
  not   g14( wr_99   ,           G176gat );
  not   g15( wr_101  ,           G204gat );
  not   g16( wr_113  ,           G64gat  );
  not   g17( wr_116  ,           G71gat  );
  not   g18( wr_118  ,           G78gat  );
  not   g19( wr_127  ,           G92gat  );
  not   g20( wr_130  ,           G99gat  );
  not   g21( wr_132  ,           G106gat );
  not   g22( wr_158  ,           G169gat );
  not   g23( wr_160  ,           G197gat );
  not   g24( wr_172  ,           G8gat   );
  not   g25( wr_175  ,           G15gat  );
  not   g26( wr_177  ,           G22gat  );
  not   g27( wr_186  ,           G36gat  );
  not   g28( wr_189  ,           G43gat  );
  not   g29( wr_191  ,           G50gat  );
  not   g30( wr_216  ,           G183gat );
  not   g31( wr_218  ,           G211gat );
  not   g32( wr_226  ,           G231gat );
  not   g33( wr_259  ,           G190gat );
  not   g34( wr_271  ,           G218gat );
  not   g35( wr_306  ,           G228gat );
  not   g36( wr_333  ,           G227gat );
  not   g37( wr_383  ,           G232gat );
  not   g38( wr_48   ,           G225gat );
  not   g39( wr_168  ,           G229gat );
  not   g40( wr_109  ,           G230gat );
  not   g41( wr_252  ,           G226gat );
  nor   g42( wr_53   , G120gat , wr_52   );
  nor   g43( wr_55   , wr_54   , G113gat );
  nor   g44( wr_58   , G134gat , wr_57   );
  nor   g45( wr_60   , wr_59   , G127gat );
  nor   g46( wr_68   , G148gat , wr_67   );
  nor   g47( wr_70   , wr_69   , G141gat );
  nor   g48( wr_73   , G162gat , wr_72   );
  nor   g49( wr_75   , wr_74   , G155gat );
  nor   g50( wr_112  , G64gat  , wr_38   );
  nor   g51( wr_114  , wr_113  , G57gat  );
  nor   g52( wr_117  , G78gat  , wr_116  );
  nor   g53( wr_119  , wr_118  , G71gat  );
  nor   g54( wr_126  , G92gat  , wr_40   );
  nor   g55( wr_128  , wr_127  , G85gat  );
  nor   g56( wr_131  , G106gat , wr_130  );
  nor   g57( wr_133  , wr_132  , G99gat  );
  nor   g58( wr_171  , G8gat   , wr_33   );
  nor   g59( wr_173  , wr_172  , G1gat   );
  nor   g60( wr_176  , G22gat  , wr_175  );
  nor   g61( wr_178  , wr_177  , G15gat  );
  nor   g62( wr_185  , G36gat  , wr_35   );
  nor   g63( wr_187  , wr_186  , G29gat  );
  nor   g64( wr_190  , G50gat  , wr_189  );
  nor   g65( wr_192  , wr_191  , G43gat  );
  nor   g66( wr_213  , G155gat , wr_57   );
  nor   g67( wr_214  , wr_72   , G127gat );
  nor   g68( wr_217  , G211gat , wr_216  );
  nor   g69( wr_219  , wr_218  , G183gat );
  nor   g70( wr_255  , G176gat , wr_158  );
  nor   g71( wr_256  , wr_99   , G169gat );
  nor   g72( wr_258  , G190gat , wr_216  );
  nor   g73( wr_260  , wr_259  , G183gat );
  nor   g74( wr_267  , G204gat , wr_160  );
  nor   g75( wr_268  , wr_101  , G197gat );
  nor   g76( wr_270  , G218gat , wr_218  );
  nor   g77( wr_272  , wr_271  , G211gat );
  nor   g78( wr_295  , G50gat  , wr_177  );
  nor   g79( wr_296  , wr_191  , G22gat  );
  nor   g80( wr_298  , G106gat , wr_118  );
  nor   g81( wr_299  , wr_132  , G78gat  );
  nor   g82( wr_322  , G43gat  , wr_175  );
  nor   g83( wr_323  , wr_189  , G15gat  );
  nor   g84( wr_325  , G99gat  , wr_116  );
  nor   g85( wr_326  , wr_130  , G71gat  );
  nor   g86( wr_372  , G162gat , wr_59   );
  nor   g87( wr_373  , wr_74   , G134gat );
  nor   g88( wr_375  , G218gat , wr_259  );
  nor   g89( wr_376  , wr_271  , G190gat );
  nor   g90( wr_227  , wr_49   , wr_226  );
  nor   g91( wr_307  , wr_49   , wr_306  );
  nor   g92( wr_334  , wr_49   , wr_333  );
  nor   g93( wr_384  , wr_49   , wr_383  );
  nor   g94( wr_34   , G29gat  , wr_33   );
  nor   g95( wr_36   , wr_35   , G1gat   );
  nor   g96( wr_39   , G85gat  , wr_38   );
  nor   g97( wr_41   , wr_40   , G57gat  );
  nor   g98( wr_155  , G141gat , wr_52   );
  nor   g99( wr_156  , wr_67   , G113gat );
  nor  g100( wr_159  , G197gat , wr_158  );
  nor  g101( wr_161  , wr_160  , G169gat );
  nor  g102( wr_50   , wr_49   , wr_48   );
  nor  g103( wr_169  , wr_49   , wr_168  );
  nor  g104( wr_96   , G148gat , wr_54   );
  nor  g105( wr_97   , wr_69   , G120gat );
  nor  g106( wr_100  , G204gat , wr_99   );
  nor  g107( wr_102  , wr_101  , G176gat );
  nor  g108( wr_241  , G36gat  , wr_172  );
  nor  g109( wr_242  , wr_186  , G8gat   );
  nor  g110( wr_244  , G92gat  , wr_113  );
  nor  g111( wr_245  , wr_127  , G64gat  );
  nor  g112( wr_110  , wr_49   , wr_109  );
  nor  g113( wr_253  , wr_49   , wr_252  );
  nor  g114( wr_56   , wr_55   , wr_53   );
  nor  g115( wr_61   , wr_60   , wr_58   );
  nor  g116( wr_71   , wr_70   , wr_68   );
  nor  g117( wr_76   , wr_75   , wr_73   );
  nor  g118( wr_115  , wr_114  , wr_112  );
  nor  g119( wr_120  , wr_119  , wr_117  );
  nor  g120( wr_129  , wr_128  , wr_126  );
  nor  g121( wr_134  , wr_133  , wr_131  );
  nor  g122( wr_174  , wr_173  , wr_171  );
  nor  g123( wr_179  , wr_178  , wr_176  );
  nor  g124( wr_188  , wr_187  , wr_185  );
  nor  g125( wr_193  , wr_192  , wr_190  );
  nor  g126( wr_257  , wr_256  , wr_255  );
  nor  g127( wr_261  , wr_260  , wr_258  );
  nor  g128( wr_269  , wr_268  , wr_267  );
  nor  g129( wr_273  , wr_272  , wr_270  );
  nor  g130( wr_215  , wr_214  , wr_213  );
  nor  g131( wr_220  , wr_219  , wr_217  );
  nor  g132( wr_297  , wr_296  , wr_295  );
  nor  g133( wr_300  , wr_299  , wr_298  );
  nor  g134( wr_324  , wr_323  , wr_322  );
  nor  g135( wr_327  , wr_326  , wr_325  );
  nor  g136( wr_374  , wr_373  , wr_372  );
  nor  g137( wr_377  , wr_376  , wr_375  );
  not  g138( wr_228  ,           wr_227  );
  not  g139( wr_308  ,           wr_307  );
  not  g140( wr_335  ,           wr_334  );
  not  g141( wr_385  ,           wr_384  );
  nor  g142( wr_37   , wr_36   , wr_34   );
  nor  g143( wr_42   , wr_41   , wr_39   );
  nor  g144( wr_157  , wr_156  , wr_155  );
  nor  g145( wr_162  , wr_161  , wr_159  );
  not  g146( wr_51   ,           wr_50   );
  not  g147( wr_170  ,           wr_169  );
  nor  g148( wr_98   , wr_97   , wr_96   );
  nor  g149( wr_103  , wr_102  , wr_100  );
  nor  g150( wr_243  , wr_242  , wr_241  );
  nor  g151( wr_246  , wr_245  , wr_244  );
  not  g152( wr_111  ,           wr_110  );
  not  g153( wr_254  ,           wr_253  );
  not  g154( wr_62   ,           wr_61   );
  not  g155( wr_64   ,           wr_56   );
  not  g156( wr_77   ,           wr_76   );
  not  g157( wr_79   ,           wr_71   );
  not  g158( wr_121  ,           wr_120  );
  not  g159( wr_123  ,           wr_115  );
  not  g160( wr_135  ,           wr_134  );
  not  g161( wr_137  ,           wr_129  );
  not  g162( wr_180  ,           wr_179  );
  not  g163( wr_182  ,           wr_174  );
  not  g164( wr_194  ,           wr_193  );
  not  g165( wr_196  ,           wr_188  );
  not  g166( wr_262  ,           wr_261  );
  not  g167( wr_264  ,           wr_257  );
  not  g168( wr_274  ,           wr_273  );
  not  g169( wr_276  ,           wr_269  );
  not  g170( wr_221  ,           wr_220  );
  not  g171( wr_223  ,           wr_215  );
  not  g172( wr_301  ,           wr_300  );
  not  g173( wr_303  ,           wr_297  );
  not  g174( wr_328  ,           wr_327  );
  not  g175( wr_330  ,           wr_324  );
  not  g176( wr_378  ,           wr_377  );
  not  g177( wr_380  ,           wr_374  );
  not  g178( wr_43   ,           wr_42   );
  not  g179( wr_45   ,           wr_37   );
  not  g180( wr_163  ,           wr_162  );
  not  g181( wr_165  ,           wr_157  );
  not  g182( wr_104  ,           wr_103  );
  not  g183( wr_106  ,           wr_98   );
  not  g184( wr_247  ,           wr_246  );
  not  g185( wr_249  ,           wr_243  );
  nor  g186( wr_63   , wr_62   , wr_56   );
  nor  g187( wr_65   , wr_61   , wr_64   );
  nor  g188( wr_78   , wr_77   , wr_71   );
  nor  g189( wr_80   , wr_76   , wr_79   );
  nor  g190( wr_122  , wr_121  , wr_115  );
  nor  g191( wr_124  , wr_120  , wr_123  );
  nor  g192( wr_136  , wr_135  , wr_129  );
  nor  g193( wr_138  , wr_134  , wr_137  );
  nor  g194( wr_181  , wr_180  , wr_174  );
  nor  g195( wr_183  , wr_179  , wr_182  );
  nor  g196( wr_195  , wr_194  , wr_188  );
  nor  g197( wr_197  , wr_193  , wr_196  );
  nor  g198( wr_263  , wr_262  , wr_257  );
  nor  g199( wr_265  , wr_261  , wr_264  );
  nor  g200( wr_275  , wr_274  , wr_269  );
  nor  g201( wr_277  , wr_273  , wr_276  );
  nor  g202( wr_222  , wr_221  , wr_215  );
  nor  g203( wr_224  , wr_220  , wr_223  );
  nor  g204( wr_302  , wr_301  , wr_297  );
  nor  g205( wr_304  , wr_300  , wr_303  );
  nor  g206( wr_329  , wr_328  , wr_324  );
  nor  g207( wr_331  , wr_327  , wr_330  );
  nor  g208( wr_379  , wr_378  , wr_374  );
  nor  g209( wr_381  , wr_377  , wr_380  );
  nor  g210( wr_44   , wr_43   , wr_37   );
  nor  g211( wr_46   , wr_42   , wr_45   );
  nor  g212( wr_164  , wr_163  , wr_157  );
  nor  g213( wr_166  , wr_162  , wr_165  );
  nor  g214( wr_105  , wr_104  , wr_98   );
  nor  g215( wr_107  , wr_103  , wr_106  );
  nor  g216( wr_248  , wr_247  , wr_243  );
  nor  g217( wr_250  , wr_246  , wr_249  );
  nor  g218( wr_66   , wr_65   , wr_63   );
  nor  g219( wr_81   , wr_80   , wr_78   );
  nor  g220( wr_125  , wr_124  , wr_122  );
  nor  g221( wr_139  , wr_138  , wr_136  );
  nor  g222( wr_184  , wr_183  , wr_181  );
  nor  g223( wr_198  , wr_197  , wr_195  );
  nor  g224( wr_266  , wr_265  , wr_263  );
  nor  g225( wr_278  , wr_277  , wr_275  );
  nor  g226( wr_225  , wr_224  , wr_222  );
  nor  g227( wr_305  , wr_304  , wr_302  );
  nor  g228( wr_332  , wr_331  , wr_329  );
  nor  g229( wr_382  , wr_381  , wr_379  );
  nor  g230( wr_47   , wr_46   , wr_44   );
  nor  g231( wr_167  , wr_166  , wr_164  );
  nor  g232( wr_108  , wr_107  , wr_105  );
  nor  g233( wr_251  , wr_250  , wr_248  );
  not  g234( wr_82   ,           wr_81   );
  not  g235( wr_84   ,           wr_66   );
  not  g236( wr_140  ,           wr_139  );
  not  g237( wr_142  ,           wr_125  );
  not  g238( wr_199  ,           wr_198  );
  not  g239( wr_201  ,           wr_184  );
  not  g240( wr_279  ,           wr_278  );
  not  g241( wr_281  ,           wr_266  );
  not  g242( wr_238  ,           wr_225  );
  not  g243( wr_318  ,           wr_305  );
  not  g244( wr_345  ,           wr_332  );
  not  g245( wr_395  ,           wr_382  );
  not  g246( wr_93   ,           wr_47   );
  not  g247( wr_210  ,           wr_167  );
  not  g248( wr_151  ,           wr_108  );
  not  g249( wr_290  ,           wr_251  );
  nor  g250( wr_229  , wr_184  , wr_142  );
  nor  g251( wr_230  , wr_201  , wr_125  );
  nor  g252( wr_309  , wr_279  , wr_81   );
  nor  g253( wr_310  , wr_278  , wr_82   );
  nor  g254( wr_336  , wr_281  , wr_66   );
  nor  g255( wr_337  , wr_266  , wr_84   );
  nor  g256( wr_386  , wr_198  , wr_140  );
  nor  g257( wr_387  , wr_199  , wr_139  );
  nor  g258( wr_83   , wr_82   , wr_66   );
  nor  g259( wr_85   , wr_81   , wr_84   );
  nor  g260( wr_200  , wr_199  , wr_184  );
  nor  g261( wr_202  , wr_198  , wr_201  );
  nor  g262( wr_141  , wr_140  , wr_125  );
  nor  g263( wr_143  , wr_139  , wr_142  );
  nor  g264( wr_280  , wr_279  , wr_266  );
  nor  g265( wr_282  , wr_278  , wr_281  );
  nor  g266( wr_231  , wr_230  , wr_229  );
  nor  g267( wr_311  , wr_310  , wr_309  );
  nor  g268( wr_338  , wr_337  , wr_336  );
  nor  g269( wr_388  , wr_387  , wr_386  );
  nor  g270( wr_86   , wr_85   , wr_83   );
  nor  g271( wr_203  , wr_202  , wr_200  );
  nor  g272( wr_144  , wr_143  , wr_141  );
  nor  g273( wr_283  , wr_282  , wr_280  );
  not  g274( wr_232  ,           wr_231  );
  not  g275( wr_312  ,           wr_311  );
  not  g276( wr_339  ,           wr_338  );
  not  g277( wr_389  ,           wr_388  );
  nor  g278( wr_234  , wr_231  , wr_227  );
  nor  g279( wr_314  , wr_311  , wr_307  );
  nor  g280( wr_341  , wr_338  , wr_334  );
  nor  g281( wr_391  , wr_388  , wr_384  );
  not  g282( wr_87   ,           wr_86   );
  not  g283( wr_204  ,           wr_203  );
  nor  g284( wr_89   , wr_86   , wr_50   );
  nor  g285( wr_206  , wr_203  , wr_169  );
  not  g286( wr_145  ,           wr_144  );
  not  g287( wr_284  ,           wr_283  );
  nor  g288( wr_147  , wr_144  , wr_110  );
  nor  g289( wr_286  , wr_283  , wr_253  );
  nor  g290( wr_233  , wr_232  , wr_228  );
  nor  g291( wr_313  , wr_312  , wr_308  );
  nor  g292( wr_340  , wr_339  , wr_335  );
  nor  g293( wr_390  , wr_389  , wr_385  );
  nor  g294( wr_88   , wr_87   , wr_51   );
  nor  g295( wr_205  , wr_204  , wr_170  );
  nor  g296( wr_146  , wr_145  , wr_111  );
  nor  g297( wr_285  , wr_284  , wr_254  );
  nor  g298( wr_235  , wr_234  , wr_233  );
  nor  g299( wr_315  , wr_314  , wr_313  );
  nor  g300( wr_342  , wr_341  , wr_340  );
  nor  g301( wr_392  , wr_391  , wr_390  );
  nor  g302( wr_90   , wr_89   , wr_88   );
  nor  g303( wr_207  , wr_206  , wr_205  );
  nor  g304( wr_148  , wr_147  , wr_146  );
  nor  g305( wr_287  , wr_286  , wr_285  );
  not  g306( wr_236  ,           wr_235  );
  not  g307( wr_316  ,           wr_315  );
  not  g308( wr_343  ,           wr_342  );
  not  g309( wr_393  ,           wr_392  );
  nor  g310( wr_239  , wr_235  , wr_238  );
  nor  g311( wr_319  , wr_315  , wr_318  );
  nor  g312( wr_346  , wr_342  , wr_345  );
  nor  g313( wr_396  , wr_392  , wr_395  );
  not  g314( wr_91   ,           wr_90   );
  not  g315( wr_208  ,           wr_207  );
  nor  g316( wr_94   , wr_90   , wr_93   );
  nor  g317( wr_211  , wr_207  , wr_210  );
  not  g318( wr_149  ,           wr_148  );
  not  g319( wr_288  ,           wr_287  );
  nor  g320( wr_152  , wr_148  , wr_151  );
  nor  g321( wr_291  , wr_287  , wr_290  );
  nor  g322( wr_237  , wr_236  , wr_225  );
  nor  g323( wr_317  , wr_316  , wr_305  );
  nor  g324( wr_344  , wr_343  , wr_332  );
  nor  g325( wr_394  , wr_393  , wr_382  );
  nor  g326( wr_92   , wr_91   , wr_47   );
  nor  g327( wr_209  , wr_208  , wr_167  );
  nor  g328( wr_150  , wr_149  , wr_108  );
  nor  g329( wr_289  , wr_288  , wr_251  );
  nor  g330( wr_240  , wr_239  , wr_237  );
  nor  g331( wr_320  , wr_319  , wr_317  );
  nor  g332( wr_347  , wr_346  , wr_344  );
  nor  g333( wr_397  , wr_396  , wr_394  );
  nor  g334( wr_95   , wr_94   , wr_92   );
  nor  g335( wr_212  , wr_211  , wr_209  );
  nor  g336( wr_153  , wr_152  , wr_150  );
  nor  g337( wr_292  , wr_291  , wr_289  );
  not  g338( wr_321  ,           wr_320  );
  not  g339( wr_353  ,           wr_347  );
  not  g340( wr_398  ,           wr_397  );
  not  g341( wr_427  ,           wr_240  );
  not  g342( wr_294  ,           wr_95   );
  not  g343( wr_456  ,           wr_212  );
  not  g344( wr_154  ,           wr_153  );
  not  g345( wr_293  ,           wr_292  );
  nor  g346( wr_359  , wr_353  , wr_321  );
  nor  g347( wr_515  , wr_398  , wr_427  );
  nor  g348( wr_354  , wr_353  , wr_320  );
  nor  g349( wr_510  , wr_397  , wr_427  );
  nor  g350( wr_348  , wr_347  , wr_321  );
  nor  g351( wr_505  , wr_398  , wr_240  );
  not  g352( wr_360  ,           wr_359  );
  not  g353( wr_516  ,           wr_515  );
  not  g354( wr_355  ,           wr_354  );
  not  g355( wr_511  ,           wr_510  );
  not  g356( wr_349  ,           wr_348  );
  not  g357( wr_506  ,           wr_505  );
  nor  g358( wr_361  , wr_360  , wr_95   );
  nor  g359( wr_364  , wr_360  , wr_294  );
  nor  g360( wr_517  , wr_516  , wr_212  );
  nor  g361( wr_520  , wr_516  , wr_456  );
  nor  g362( wr_356  , wr_355  , wr_294  );
  nor  g363( wr_512  , wr_511  , wr_456  );
  nor  g364( wr_350  , wr_349  , wr_294  );
  nor  g365( wr_507  , wr_506  , wr_456  );
  not  g366( wr_362  ,           wr_361  );
  not  g367( wr_365  ,           wr_364  );
  not  g368( wr_518  ,           wr_517  );
  not  g369( wr_521  ,           wr_520  );
  not  g370( wr_357  ,           wr_356  );
  not  g371( wr_513  ,           wr_512  );
  not  g372( wr_351  ,           wr_350  );
  not  g373( wr_508  ,           wr_507  );
  nor  g374( wr_363  , wr_362  , wr_293  );
  nor  g375( wr_366  , wr_365  , wr_292  );
  nor  g376( wr_519  , wr_518  , wr_154  );
  nor  g377( wr_522  , wr_521  , wr_153  );
  nor  g378( wr_358  , wr_357  , wr_293  );
  nor  g379( wr_514  , wr_513  , wr_154  );
  nor  g380( wr_352  , wr_351  , wr_293  );
  nor  g381( wr_509  , wr_508  , wr_154  );
  nor  g382( wr_367  , wr_366  , wr_363  );
  nor  g383( wr_523  , wr_522  , wr_519  );
  not  g384( wr_368  ,           wr_367  );
  not  g385( wr_524  ,           wr_523  );
  nor  g386( wr_369  , wr_368  , wr_358  );
  nor  g387( wr_525  , wr_524  , wr_514  );
  not  g388( wr_370  ,           wr_369  );
  not  g389( wr_526  ,           wr_525  );
  nor  g390( wr_371  , wr_370  , wr_352  );
  nor  g391( wr_527  , wr_526  , wr_509  );
  nor  g392( wr_399  , wr_398  , wr_371  );
  nor  g393( wr_428  , wr_397  , wr_371  );
  nor  g394( wr_528  , wr_527  , wr_321  );
  nor  g395( wr_556  , wr_527  , wr_320  );
  not  g396( wr_400  ,           wr_399  );
  not  g397( wr_429  ,           wr_428  );
  not  g398( wr_529  ,           wr_528  );
  not  g399( wr_557  ,           wr_556  );
  nor  g400( wr_401  , wr_400  , wr_240  );
  nor  g401( wr_430  , wr_429  , wr_427  );
  nor  g402( wr_530  , wr_529  , wr_347  );
  nor  g403( wr_558  , wr_557  , wr_353  );
  not  g404( wr_402  ,           wr_401  );
  not  g405( wr_431  ,           wr_430  );
  not  g406( wr_531  ,           wr_530  );
  not  g407( wr_559  ,           wr_558  );
  nor  g408( wr_403  , wr_402  , wr_212  );
  nor  g409( wr_432  , wr_431  , wr_212  );
  nor  g410( wr_457  , wr_402  , wr_456  );
  nor  g411( wr_481  , wr_431  , wr_456  );
  nor  g412( wr_532  , wr_531  , wr_95   );
  nor  g413( wr_560  , wr_559  , wr_95   );
  nor  g414( wr_584  , wr_531  , wr_294  );
  nor  g415( wr_608  , wr_559  , wr_294  );
  not  g416( wr_404  ,           wr_403  );
  not  g417( wr_433  ,           wr_432  );
  not  g418( wr_458  ,           wr_457  );
  not  g419( wr_482  ,           wr_481  );
  not  g420( wr_533  ,           wr_532  );
  not  g421( wr_561  ,           wr_560  );
  not  g422( wr_585  ,           wr_584  );
  not  g423( wr_609  ,           wr_608  );
  nor  g424( wr_405  , wr_404  , wr_154  );
  nor  g425( wr_434  , wr_433  , wr_154  );
  nor  g426( wr_459  , wr_458  , wr_153  );
  nor  g427( wr_483  , wr_482  , wr_153  );
  nor  g428( wr_534  , wr_533  , wr_293  );
  nor  g429( wr_562  , wr_561  , wr_293  );
  nor  g430( wr_586  , wr_585  , wr_292  );
  nor  g431( wr_610  , wr_609  , wr_292  );
  not  g432( wr_406  ,           wr_405  );
  not  g433( wr_435  ,           wr_434  );
  not  g434( wr_460  ,           wr_459  );
  not  g435( wr_484  ,           wr_483  );
  not  g436( wr_535  ,           wr_534  );
  not  g437( wr_563  ,           wr_562  );
  not  g438( wr_587  ,           wr_586  );
  not  g439( wr_611  ,           wr_610  );
  nor  g440( wr_407  , wr_406  , wr_95   );
  nor  g441( wr_412  , wr_406  , wr_292  );
  nor  g442( wr_417  , wr_406  , wr_347  );
  nor  g443( wr_422  , wr_406  , wr_320  );
  nor  g444( wr_436  , wr_435  , wr_95   );
  nor  g445( wr_441  , wr_435  , wr_292  );
  nor  g446( wr_446  , wr_435  , wr_347  );
  nor  g447( wr_451  , wr_435  , wr_320  );
  nor  g448( wr_461  , wr_460  , wr_95   );
  nor  g449( wr_466  , wr_460  , wr_292  );
  nor  g450( wr_471  , wr_460  , wr_347  );
  nor  g451( wr_476  , wr_460  , wr_320  );
  nor  g452( wr_485  , wr_484  , wr_95   );
  nor  g453( wr_490  , wr_484  , wr_292  );
  nor  g454( wr_495  , wr_484  , wr_347  );
  nor  g455( wr_500  , wr_484  , wr_320  );
  nor  g456( wr_536  , wr_535  , wr_212  );
  nor  g457( wr_541  , wr_535  , wr_153  );
  nor  g458( wr_546  , wr_535  , wr_240  );
  nor  g459( wr_551  , wr_535  , wr_397  );
  nor  g460( wr_564  , wr_563  , wr_212  );
  nor  g461( wr_569  , wr_563  , wr_153  );
  nor  g462( wr_574  , wr_563  , wr_240  );
  nor  g463( wr_579  , wr_563  , wr_397  );
  nor  g464( wr_588  , wr_587  , wr_212  );
  nor  g465( wr_593  , wr_587  , wr_153  );
  nor  g466( wr_598  , wr_587  , wr_240  );
  nor  g467( wr_603  , wr_587  , wr_397  );
  nor  g468( wr_612  , wr_611  , wr_212  );
  nor  g469( wr_617  , wr_611  , wr_153  );
  nor  g470( wr_622  , wr_611  , wr_240  );
  nor  g471( wr_627  , wr_611  , wr_397  );
  not  g472( wr_409  ,           wr_407  );
  not  g473( wr_414  ,           wr_412  );
  not  g474( wr_419  ,           wr_417  );
  not  g475( wr_424  ,           wr_422  );
  not  g476( wr_438  ,           wr_436  );
  not  g477( wr_443  ,           wr_441  );
  not  g478( wr_448  ,           wr_446  );
  not  g479( wr_453  ,           wr_451  );
  not  g480( wr_463  ,           wr_461  );
  not  g481( wr_468  ,           wr_466  );
  not  g482( wr_473  ,           wr_471  );
  not  g483( wr_478  ,           wr_476  );
  not  g484( wr_487  ,           wr_485  );
  not  g485( wr_492  ,           wr_490  );
  not  g486( wr_497  ,           wr_495  );
  not  g487( wr_502  ,           wr_500  );
  not  g488( wr_538  ,           wr_536  );
  not  g489( wr_543  ,           wr_541  );
  not  g490( wr_548  ,           wr_546  );
  not  g491( wr_553  ,           wr_551  );
  not  g492( wr_566  ,           wr_564  );
  not  g493( wr_571  ,           wr_569  );
  not  g494( wr_576  ,           wr_574  );
  not  g495( wr_581  ,           wr_579  );
  not  g496( wr_590  ,           wr_588  );
  not  g497( wr_595  ,           wr_593  );
  not  g498( wr_600  ,           wr_598  );
  not  g499( wr_605  ,           wr_603  );
  not  g500( wr_614  ,           wr_612  );
  not  g501( wr_619  ,           wr_617  );
  not  g502( wr_624  ,           wr_622  );
  not  g503( wr_629  ,           wr_627  );
  nor  g504( wr_408  , wr_407  , wr_33   );
  nor  g505( wr_413  , wr_412  , wr_172  );
  nor  g506( wr_418  , wr_417  , wr_175  );
  nor  g507( wr_423  , wr_422  , wr_177  );
  nor  g508( wr_437  , wr_436  , wr_35   );
  nor  g509( wr_442  , wr_441  , wr_186  );
  nor  g510( wr_447  , wr_446  , wr_189  );
  nor  g511( wr_452  , wr_451  , wr_191  );
  nor  g512( wr_462  , wr_461  , wr_38   );
  nor  g513( wr_467  , wr_466  , wr_113  );
  nor  g514( wr_472  , wr_471  , wr_116  );
  nor  g515( wr_477  , wr_476  , wr_118  );
  nor  g516( wr_486  , wr_485  , wr_40   );
  nor  g517( wr_491  , wr_490  , wr_127  );
  nor  g518( wr_496  , wr_495  , wr_130  );
  nor  g519( wr_501  , wr_500  , wr_132  );
  nor  g520( wr_537  , wr_536  , wr_52   );
  nor  g521( wr_542  , wr_541  , wr_54   );
  nor  g522( wr_547  , wr_546  , wr_57   );
  nor  g523( wr_552  , wr_551  , wr_59   );
  nor  g524( wr_565  , wr_564  , wr_67   );
  nor  g525( wr_570  , wr_569  , wr_69   );
  nor  g526( wr_575  , wr_574  , wr_72   );
  nor  g527( wr_580  , wr_579  , wr_74   );
  nor  g528( wr_589  , wr_588  , wr_158  );
  nor  g529( wr_594  , wr_593  , wr_99   );
  nor  g530( wr_599  , wr_598  , wr_216  );
  nor  g531( wr_604  , wr_603  , wr_259  );
  nor  g532( wr_613  , wr_612  , wr_160  );
  nor  g533( wr_618  , wr_617  , wr_101  );
  nor  g534( wr_623  , wr_622  , wr_218  );
  nor  g535( wr_628  , wr_627  , wr_271  );
  nor  g536( wr_410  , wr_409  , G1gat   );
  nor  g537( wr_415  , wr_414  , G8gat   );
  nor  g538( wr_420  , wr_419  , G15gat  );
  nor  g539( wr_425  , wr_424  , G22gat  );
  nor  g540( wr_439  , wr_438  , G29gat  );
  nor  g541( wr_444  , wr_443  , G36gat  );
  nor  g542( wr_449  , wr_448  , G43gat  );
  nor  g543( wr_454  , wr_453  , G50gat  );
  nor  g544( wr_464  , wr_463  , G57gat  );
  nor  g545( wr_469  , wr_468  , G64gat  );
  nor  g546( wr_474  , wr_473  , G71gat  );
  nor  g547( wr_479  , wr_478  , G78gat  );
  nor  g548( wr_488  , wr_487  , G85gat  );
  nor  g549( wr_493  , wr_492  , G92gat  );
  nor  g550( wr_498  , wr_497  , G99gat  );
  nor  g551( wr_503  , wr_502  , G106gat );
  nor  g552( wr_539  , wr_538  , G113gat );
  nor  g553( wr_544  , wr_543  , G120gat );
  nor  g554( wr_549  , wr_548  , G127gat );
  nor  g555( wr_554  , wr_553  , G134gat );
  nor  g556( wr_567  , wr_566  , G141gat );
  nor  g557( wr_572  , wr_571  , G148gat );
  nor  g558( wr_577  , wr_576  , G155gat );
  nor  g559( wr_582  , wr_581  , G162gat );
  nor  g560( wr_591  , wr_590  , G169gat );
  nor  g561( wr_596  , wr_595  , G176gat );
  nor  g562( wr_601  , wr_600  , G183gat );
  nor  g563( wr_606  , wr_605  , G190gat );
  nor  g564( wr_615  , wr_614  , G197gat );
  nor  g565( wr_620  , wr_619  , G204gat );
  nor  g566( wr_625  , wr_624  , G211gat );
  nor  g567( wr_630  , wr_629  , G218gat );
  nor  g568( wr_411  , wr_410  , wr_408  );
  nor  g569( wr_416  , wr_415  , wr_413  );
  nor  g570( wr_421  , wr_420  , wr_418  );
  nor  g571( wr_426  , wr_425  , wr_423  );
  nor  g572( wr_440  , wr_439  , wr_437  );
  nor  g573( wr_445  , wr_444  , wr_442  );
  nor  g574( wr_450  , wr_449  , wr_447  );
  nor  g575( wr_455  , wr_454  , wr_452  );
  nor  g576( wr_465  , wr_464  , wr_462  );
  nor  g577( wr_470  , wr_469  , wr_467  );
  nor  g578( wr_475  , wr_474  , wr_472  );
  nor  g579( wr_480  , wr_479  , wr_477  );
  nor  g580( wr_489  , wr_488  , wr_486  );
  nor  g581( wr_494  , wr_493  , wr_491  );
  nor  g582( wr_499  , wr_498  , wr_496  );
  nor  g583( wr_504  , wr_503  , wr_501  );
  nor  g584( wr_540  , wr_539  , wr_537  );
  nor  g585( wr_545  , wr_544  , wr_542  );
  nor  g586( wr_550  , wr_549  , wr_547  );
  nor  g587( wr_555  , wr_554  , wr_552  );
  nor  g588( wr_568  , wr_567  , wr_565  );
  nor  g589( wr_573  , wr_572  , wr_570  );
  nor  g590( wr_578  , wr_577  , wr_575  );
  nor  g591( wr_583  , wr_582  , wr_580  );
  nor  g592( wr_592  , wr_591  , wr_589  );
  nor  g593( wr_597  , wr_596  , wr_594  );
  nor  g594( wr_602  , wr_601  , wr_599  );
  nor  g595( wr_607  , wr_606  , wr_604  );
  nor  g596( wr_616  , wr_615  , wr_613  );
  nor  g597( wr_621  , wr_620  , wr_618  );
  nor  g598( wr_626  , wr_625  , wr_623  );
  nor  g599( wr_631  , wr_630  , wr_628  );
  not  g600( G1324gat,           wr_411  );
  not  g601( G1325gat,           wr_416  );
  not  g602( G1326gat,           wr_421  );
  not  g603( G1327gat,           wr_426  );
  not  g604( G1328gat,           wr_440  );
  not  g605( G1329gat,           wr_445  );
  not  g606( G1330gat,           wr_450  );
  not  g607( G1331gat,           wr_455  );
  not  g608( G1332gat,           wr_465  );
  not  g609( G1333gat,           wr_470  );
  not  g610( G1334gat,           wr_475  );
  not  g611( G1335gat,           wr_480  );
  not  g612( G1336gat,           wr_489  );
  not  g613( G1337gat,           wr_494  );
  not  g614( G1338gat,           wr_499  );
  not  g615( G1339gat,           wr_504  );
  not  g616( G1340gat,           wr_540  );
  not  g617( G1341gat,           wr_545  );
  not  g618( G1342gat,           wr_550  );
  not  g619( G1343gat,           wr_555  );
  not  g620( G1344gat,           wr_568  );
  not  g621( G1345gat,           wr_573  );
  not  g622( G1346gat,           wr_578  );
  not  g623( G1347gat,           wr_583  );
  not  g624( G1348gat,           wr_592  );
  not  g625( G1349gat,           wr_597  );
  not  g626( G1350gat,           wr_602  );
  not  g627( G1351gat,           wr_607  );
  not  g628( G1352gat,           wr_616  );
  not  g629( G1353gat,           wr_621  );
  not  g630( G1354gat,           wr_626  );
  not  g631( G1355gat,           wr_631  );

endmodule
